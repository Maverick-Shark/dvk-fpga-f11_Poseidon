
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"aa",x"b7",x"c0",x"4a"),
     1 => (x"c2",x"87",x"d3",x"03"),
     2 => (x"05",x"bf",x"cd",x"cd"),
     3 => (x"4b",x"c1",x"87",x"c4"),
     4 => (x"4b",x"c0",x"87",x"c2"),
     5 => (x"5b",x"d1",x"cd",x"c2"),
     6 => (x"cd",x"c2",x"87",x"c4"),
     7 => (x"cd",x"c2",x"5a",x"d1"),
     8 => (x"c1",x"4a",x"bf",x"cd"),
     9 => (x"a2",x"c0",x"c1",x"9a"),
    10 => (x"87",x"e8",x"ec",x"49"),
    11 => (x"cd",x"c2",x"48",x"fc"),
    12 => (x"fe",x"78",x"bf",x"cd"),
    13 => (x"71",x"1e",x"87",x"ef"),
    14 => (x"1e",x"66",x"c4",x"4a"),
    15 => (x"fd",x"e9",x"49",x"72"),
    16 => (x"4f",x"26",x"26",x"87"),
    17 => (x"cd",x"cd",x"c2",x"1e"),
    18 => (x"d7",x"e6",x"49",x"bf"),
    19 => (x"d6",x"ec",x"c2",x"87"),
    20 => (x"78",x"bf",x"e8",x"48"),
    21 => (x"48",x"d2",x"ec",x"c2"),
    22 => (x"c2",x"78",x"bf",x"ec"),
    23 => (x"4a",x"bf",x"d6",x"ec"),
    24 => (x"99",x"ff",x"c3",x"49"),
    25 => (x"72",x"2a",x"b7",x"c8"),
    26 => (x"c2",x"b0",x"71",x"48"),
    27 => (x"26",x"58",x"de",x"ec"),
    28 => (x"5b",x"5e",x"0e",x"4f"),
    29 => (x"71",x"0e",x"5d",x"5c"),
    30 => (x"87",x"c8",x"ff",x"4b"),
    31 => (x"48",x"d1",x"ec",x"c2"),
    32 => (x"49",x"73",x"50",x"c0"),
    33 => (x"70",x"87",x"fd",x"e5"),
    34 => (x"9c",x"c2",x"4c",x"49"),
    35 => (x"cb",x"49",x"ee",x"cb"),
    36 => (x"49",x"70",x"87",x"c3"),
    37 => (x"d1",x"ec",x"c2",x"4d"),
    38 => (x"c1",x"05",x"bf",x"97"),
    39 => (x"66",x"d0",x"87",x"e2"),
    40 => (x"da",x"ec",x"c2",x"49"),
    41 => (x"d6",x"05",x"99",x"bf"),
    42 => (x"49",x"66",x"d4",x"87"),
    43 => (x"bf",x"d2",x"ec",x"c2"),
    44 => (x"87",x"cb",x"05",x"99"),
    45 => (x"cb",x"e5",x"49",x"73"),
    46 => (x"02",x"98",x"70",x"87"),
    47 => (x"c1",x"87",x"c1",x"c1"),
    48 => (x"87",x"c0",x"fe",x"4c"),
    49 => (x"d8",x"ca",x"49",x"75"),
    50 => (x"02",x"98",x"70",x"87"),
    51 => (x"ec",x"c2",x"87",x"c6"),
    52 => (x"50",x"c1",x"48",x"d1"),
    53 => (x"97",x"d1",x"ec",x"c2"),
    54 => (x"e3",x"c0",x"05",x"bf"),
    55 => (x"da",x"ec",x"c2",x"87"),
    56 => (x"66",x"d0",x"49",x"bf"),
    57 => (x"d6",x"ff",x"05",x"99"),
    58 => (x"d2",x"ec",x"c2",x"87"),
    59 => (x"66",x"d4",x"49",x"bf"),
    60 => (x"ca",x"ff",x"05",x"99"),
    61 => (x"e4",x"49",x"73",x"87"),
    62 => (x"98",x"70",x"87",x"ca"),
    63 => (x"87",x"ff",x"fe",x"05"),
    64 => (x"dc",x"fb",x"48",x"74"),
    65 => (x"5b",x"5e",x"0e",x"87"),
    66 => (x"f4",x"0e",x"5d",x"5c"),
    67 => (x"4c",x"4d",x"c0",x"86"),
    68 => (x"c4",x"7e",x"bf",x"ec"),
    69 => (x"ec",x"c2",x"48",x"a6"),
    70 => (x"c1",x"78",x"bf",x"de"),
    71 => (x"c7",x"1e",x"c0",x"1e"),
    72 => (x"87",x"cd",x"fd",x"49"),
    73 => (x"98",x"70",x"86",x"c8"),
    74 => (x"ff",x"87",x"cd",x"02"),
    75 => (x"87",x"cc",x"fb",x"49"),
    76 => (x"e3",x"49",x"da",x"c1"),
    77 => (x"4d",x"c1",x"87",x"ce"),
    78 => (x"97",x"d1",x"ec",x"c2"),
    79 => (x"87",x"c3",x"02",x"bf"),
    80 => (x"c2",x"87",x"fe",x"d4"),
    81 => (x"4b",x"bf",x"d6",x"ec"),
    82 => (x"bf",x"cd",x"cd",x"c2"),
    83 => (x"87",x"e9",x"c0",x"05"),
    84 => (x"e2",x"49",x"fd",x"c3"),
    85 => (x"fa",x"c3",x"87",x"ee"),
    86 => (x"87",x"e8",x"e2",x"49"),
    87 => (x"ff",x"c3",x"49",x"73"),
    88 => (x"c0",x"1e",x"71",x"99"),
    89 => (x"87",x"ce",x"fb",x"49"),
    90 => (x"b7",x"c8",x"49",x"73"),
    91 => (x"c1",x"1e",x"71",x"29"),
    92 => (x"87",x"c2",x"fb",x"49"),
    93 => (x"fa",x"c5",x"86",x"c8"),
    94 => (x"da",x"ec",x"c2",x"87"),
    95 => (x"02",x"9b",x"4b",x"bf"),
    96 => (x"cd",x"c2",x"87",x"dd"),
    97 => (x"c7",x"49",x"bf",x"c9"),
    98 => (x"98",x"70",x"87",x"d7"),
    99 => (x"c0",x"87",x"c4",x"05"),
   100 => (x"c2",x"87",x"d2",x"4b"),
   101 => (x"fc",x"c6",x"49",x"e0"),
   102 => (x"cd",x"cd",x"c2",x"87"),
   103 => (x"c2",x"87",x"c6",x"58"),
   104 => (x"c0",x"48",x"c9",x"cd"),
   105 => (x"c2",x"49",x"73",x"78"),
   106 => (x"87",x"cd",x"05",x"99"),
   107 => (x"e1",x"49",x"eb",x"c3"),
   108 => (x"49",x"70",x"87",x"d2"),
   109 => (x"c2",x"02",x"99",x"c2"),
   110 => (x"73",x"4c",x"fb",x"87"),
   111 => (x"05",x"99",x"c1",x"49"),
   112 => (x"f4",x"c3",x"87",x"cd"),
   113 => (x"87",x"fc",x"e0",x"49"),
   114 => (x"99",x"c2",x"49",x"70"),
   115 => (x"fa",x"87",x"c2",x"02"),
   116 => (x"c8",x"49",x"73",x"4c"),
   117 => (x"87",x"cd",x"05",x"99"),
   118 => (x"e0",x"49",x"f5",x"c3"),
   119 => (x"49",x"70",x"87",x"e6"),
   120 => (x"d4",x"02",x"99",x"c2"),
   121 => (x"e2",x"ec",x"c2",x"87"),
   122 => (x"87",x"c9",x"02",x"bf"),
   123 => (x"c2",x"88",x"c1",x"48"),
   124 => (x"c2",x"58",x"e6",x"ec"),
   125 => (x"c1",x"4c",x"ff",x"87"),
   126 => (x"c4",x"49",x"73",x"4d"),
   127 => (x"87",x"ce",x"05",x"99"),
   128 => (x"ff",x"49",x"f2",x"c3"),
   129 => (x"70",x"87",x"fd",x"df"),
   130 => (x"02",x"99",x"c2",x"49"),
   131 => (x"ec",x"c2",x"87",x"db"),
   132 => (x"48",x"7e",x"bf",x"e2"),
   133 => (x"03",x"a8",x"b7",x"c7"),
   134 => (x"48",x"6e",x"87",x"cb"),
   135 => (x"ec",x"c2",x"80",x"c1"),
   136 => (x"c2",x"c0",x"58",x"e6"),
   137 => (x"c1",x"4c",x"fe",x"87"),
   138 => (x"49",x"fd",x"c3",x"4d"),
   139 => (x"87",x"d4",x"df",x"ff"),
   140 => (x"99",x"c2",x"49",x"70"),
   141 => (x"c2",x"87",x"d5",x"02"),
   142 => (x"02",x"bf",x"e2",x"ec"),
   143 => (x"c2",x"87",x"c9",x"c0"),
   144 => (x"c0",x"48",x"e2",x"ec"),
   145 => (x"87",x"c2",x"c0",x"78"),
   146 => (x"4d",x"c1",x"4c",x"fd"),
   147 => (x"ff",x"49",x"fa",x"c3"),
   148 => (x"70",x"87",x"f1",x"de"),
   149 => (x"02",x"99",x"c2",x"49"),
   150 => (x"ec",x"c2",x"87",x"d9"),
   151 => (x"c7",x"48",x"bf",x"e2"),
   152 => (x"c0",x"03",x"a8",x"b7"),
   153 => (x"ec",x"c2",x"87",x"c9"),
   154 => (x"78",x"c7",x"48",x"e2"),
   155 => (x"fc",x"87",x"c2",x"c0"),
   156 => (x"c0",x"4d",x"c1",x"4c"),
   157 => (x"c0",x"03",x"ac",x"b7"),
   158 => (x"66",x"c4",x"87",x"d1"),
   159 => (x"82",x"d8",x"c1",x"4a"),
   160 => (x"c6",x"c0",x"02",x"6a"),
   161 => (x"74",x"4b",x"6a",x"87"),
   162 => (x"c0",x"0f",x"73",x"49"),
   163 => (x"1e",x"f0",x"c3",x"1e"),
   164 => (x"f7",x"49",x"da",x"c1"),
   165 => (x"86",x"c8",x"87",x"db"),
   166 => (x"c0",x"02",x"98",x"70"),
   167 => (x"a6",x"c8",x"87",x"e2"),
   168 => (x"e2",x"ec",x"c2",x"48"),
   169 => (x"66",x"c8",x"78",x"bf"),
   170 => (x"c4",x"91",x"cb",x"49"),
   171 => (x"80",x"71",x"48",x"66"),
   172 => (x"bf",x"6e",x"7e",x"70"),
   173 => (x"87",x"c8",x"c0",x"02"),
   174 => (x"c8",x"4b",x"bf",x"6e"),
   175 => (x"0f",x"73",x"49",x"66"),
   176 => (x"c0",x"02",x"9d",x"75"),
   177 => (x"ec",x"c2",x"87",x"c8"),
   178 => (x"f3",x"49",x"bf",x"e2"),
   179 => (x"cd",x"c2",x"87",x"c9"),
   180 => (x"c0",x"02",x"bf",x"d1"),
   181 => (x"c2",x"49",x"87",x"dd"),
   182 => (x"98",x"70",x"87",x"c7"),
   183 => (x"87",x"d3",x"c0",x"02"),
   184 => (x"bf",x"e2",x"ec",x"c2"),
   185 => (x"87",x"ef",x"f2",x"49"),
   186 => (x"cf",x"f4",x"49",x"c0"),
   187 => (x"d1",x"cd",x"c2",x"87"),
   188 => (x"f4",x"78",x"c0",x"48"),
   189 => (x"87",x"e9",x"f3",x"8e"),
   190 => (x"5c",x"5b",x"5e",x"0e"),
   191 => (x"71",x"1e",x"0e",x"5d"),
   192 => (x"de",x"ec",x"c2",x"4c"),
   193 => (x"cd",x"c1",x"49",x"bf"),
   194 => (x"d1",x"c1",x"4d",x"a1"),
   195 => (x"74",x"7e",x"69",x"81"),
   196 => (x"87",x"cf",x"02",x"9c"),
   197 => (x"74",x"4b",x"a5",x"c4"),
   198 => (x"de",x"ec",x"c2",x"7b"),
   199 => (x"c8",x"f3",x"49",x"bf"),
   200 => (x"74",x"7b",x"6e",x"87"),
   201 => (x"87",x"c4",x"05",x"9c"),
   202 => (x"87",x"c2",x"4b",x"c0"),
   203 => (x"49",x"73",x"4b",x"c1"),
   204 => (x"d4",x"87",x"c9",x"f3"),
   205 => (x"87",x"c7",x"02",x"66"),
   206 => (x"70",x"87",x"da",x"49"),
   207 => (x"c0",x"87",x"c2",x"4a"),
   208 => (x"d5",x"cd",x"c2",x"4a"),
   209 => (x"d8",x"f2",x"26",x"5a"),
   210 => (x"00",x"00",x"00",x"87"),
   211 => (x"00",x"00",x"00",x"00"),
   212 => (x"00",x"00",x"00",x"00"),
   213 => (x"4a",x"71",x"1e",x"00"),
   214 => (x"49",x"bf",x"c8",x"ff"),
   215 => (x"26",x"48",x"a1",x"72"),
   216 => (x"c8",x"ff",x"1e",x"4f"),
   217 => (x"c0",x"fe",x"89",x"bf"),
   218 => (x"c0",x"c0",x"c0",x"c0"),
   219 => (x"87",x"c4",x"01",x"a9"),
   220 => (x"87",x"c2",x"4a",x"c0"),
   221 => (x"48",x"72",x"4a",x"c1"),
   222 => (x"5e",x"0e",x"4f",x"26"),
   223 => (x"0e",x"5d",x"5c",x"5b"),
   224 => (x"d4",x"ff",x"4b",x"71"),
   225 => (x"48",x"66",x"d0",x"4c"),
   226 => (x"49",x"d6",x"78",x"c0"),
   227 => (x"87",x"f4",x"db",x"ff"),
   228 => (x"6c",x"7c",x"ff",x"c3"),
   229 => (x"99",x"ff",x"c3",x"49"),
   230 => (x"c3",x"49",x"4d",x"71"),
   231 => (x"e0",x"c1",x"99",x"f0"),
   232 => (x"87",x"cb",x"05",x"a9"),
   233 => (x"6c",x"7c",x"ff",x"c3"),
   234 => (x"d0",x"98",x"c3",x"48"),
   235 => (x"c3",x"78",x"08",x"66"),
   236 => (x"4a",x"6c",x"7c",x"ff"),
   237 => (x"c3",x"31",x"c8",x"49"),
   238 => (x"4a",x"6c",x"7c",x"ff"),
   239 => (x"49",x"72",x"b2",x"71"),
   240 => (x"ff",x"c3",x"31",x"c8"),
   241 => (x"71",x"4a",x"6c",x"7c"),
   242 => (x"c8",x"49",x"72",x"b2"),
   243 => (x"7c",x"ff",x"c3",x"31"),
   244 => (x"b2",x"71",x"4a",x"6c"),
   245 => (x"c0",x"48",x"d0",x"ff"),
   246 => (x"9b",x"73",x"78",x"e0"),
   247 => (x"72",x"87",x"c2",x"02"),
   248 => (x"26",x"48",x"75",x"7b"),
   249 => (x"26",x"4c",x"26",x"4d"),
   250 => (x"1e",x"4f",x"26",x"4b"),
   251 => (x"5e",x"0e",x"4f",x"26"),
   252 => (x"f8",x"0e",x"5c",x"5b"),
   253 => (x"c8",x"1e",x"76",x"86"),
   254 => (x"fd",x"fd",x"49",x"a6"),
   255 => (x"70",x"86",x"c4",x"87"),
   256 => (x"c0",x"48",x"6e",x"4b"),
   257 => (x"c6",x"c3",x"01",x"a8"),
   258 => (x"c3",x"4a",x"73",x"87"),
   259 => (x"d0",x"c1",x"9a",x"f0"),
   260 => (x"87",x"c7",x"02",x"aa"),
   261 => (x"05",x"aa",x"e0",x"c1"),
   262 => (x"73",x"87",x"f4",x"c2"),
   263 => (x"02",x"99",x"c8",x"49"),
   264 => (x"c6",x"ff",x"87",x"c3"),
   265 => (x"c3",x"4c",x"73",x"87"),
   266 => (x"05",x"ac",x"c2",x"9c"),
   267 => (x"c4",x"87",x"cd",x"c1"),
   268 => (x"31",x"c9",x"49",x"66"),
   269 => (x"66",x"c4",x"1e",x"71"),
   270 => (x"c2",x"92",x"d4",x"4a"),
   271 => (x"72",x"49",x"e6",x"ec"),
   272 => (x"e0",x"d5",x"fe",x"81"),
   273 => (x"49",x"66",x"c4",x"87"),
   274 => (x"49",x"e3",x"c0",x"1e"),
   275 => (x"87",x"d9",x"d9",x"ff"),
   276 => (x"d8",x"ff",x"49",x"d8"),
   277 => (x"c0",x"c8",x"87",x"ee"),
   278 => (x"d6",x"db",x"c2",x"1e"),
   279 => (x"f5",x"f1",x"fd",x"49"),
   280 => (x"48",x"d0",x"ff",x"87"),
   281 => (x"c2",x"78",x"e0",x"c0"),
   282 => (x"d0",x"1e",x"d6",x"db"),
   283 => (x"92",x"d4",x"4a",x"66"),
   284 => (x"49",x"e6",x"ec",x"c2"),
   285 => (x"d3",x"fe",x"81",x"72"),
   286 => (x"86",x"d0",x"87",x"e8"),
   287 => (x"c1",x"05",x"ac",x"c1"),
   288 => (x"66",x"c4",x"87",x"cd"),
   289 => (x"71",x"31",x"c9",x"49"),
   290 => (x"4a",x"66",x"c4",x"1e"),
   291 => (x"ec",x"c2",x"92",x"d4"),
   292 => (x"81",x"72",x"49",x"e6"),
   293 => (x"87",x"cd",x"d4",x"fe"),
   294 => (x"1e",x"d6",x"db",x"c2"),
   295 => (x"d4",x"4a",x"66",x"c8"),
   296 => (x"e6",x"ec",x"c2",x"92"),
   297 => (x"fe",x"81",x"72",x"49"),
   298 => (x"c8",x"87",x"f4",x"d1"),
   299 => (x"c0",x"1e",x"49",x"66"),
   300 => (x"d7",x"ff",x"49",x"e3"),
   301 => (x"49",x"d7",x"87",x"f3"),
   302 => (x"87",x"c8",x"d7",x"ff"),
   303 => (x"c2",x"1e",x"c0",x"c8"),
   304 => (x"fd",x"49",x"d6",x"db"),
   305 => (x"d0",x"87",x"fe",x"ef"),
   306 => (x"48",x"d0",x"ff",x"86"),
   307 => (x"f8",x"78",x"e0",x"c0"),
   308 => (x"87",x"d1",x"fc",x"8e"),
   309 => (x"5c",x"5b",x"5e",x"0e"),
   310 => (x"71",x"1e",x"0e",x"5d"),
   311 => (x"4c",x"d4",x"ff",x"4d"),
   312 => (x"48",x"7e",x"66",x"d4"),
   313 => (x"06",x"a8",x"b7",x"c3"),
   314 => (x"48",x"c0",x"87",x"c5"),
   315 => (x"75",x"87",x"e2",x"c1"),
   316 => (x"c1",x"e2",x"fe",x"49"),
   317 => (x"c4",x"1e",x"75",x"87"),
   318 => (x"93",x"d4",x"4b",x"66"),
   319 => (x"83",x"e6",x"ec",x"c2"),
   320 => (x"cc",x"fe",x"49",x"73"),
   321 => (x"83",x"c8",x"87",x"fd"),
   322 => (x"d0",x"ff",x"4b",x"6b"),
   323 => (x"78",x"e1",x"c8",x"48"),
   324 => (x"49",x"73",x"7c",x"dd"),
   325 => (x"71",x"99",x"ff",x"c3"),
   326 => (x"c8",x"49",x"73",x"7c"),
   327 => (x"ff",x"c3",x"29",x"b7"),
   328 => (x"73",x"7c",x"71",x"99"),
   329 => (x"29",x"b7",x"d0",x"49"),
   330 => (x"71",x"99",x"ff",x"c3"),
   331 => (x"d8",x"49",x"73",x"7c"),
   332 => (x"7c",x"71",x"29",x"b7"),
   333 => (x"7c",x"7c",x"7c",x"c0"),
   334 => (x"7c",x"7c",x"7c",x"7c"),
   335 => (x"7c",x"7c",x"7c",x"7c"),
   336 => (x"78",x"e0",x"c0",x"7c"),
   337 => (x"dc",x"1e",x"66",x"c4"),
   338 => (x"dc",x"d5",x"ff",x"49"),
   339 => (x"73",x"86",x"c8",x"87"),
   340 => (x"ce",x"fa",x"26",x"48"),
   341 => (x"5b",x"5e",x"0e",x"87"),
   342 => (x"1e",x"0e",x"5d",x"5c"),
   343 => (x"d4",x"ff",x"7e",x"71"),
   344 => (x"c2",x"1e",x"6e",x"4b"),
   345 => (x"fe",x"49",x"fa",x"ec"),
   346 => (x"c4",x"87",x"d8",x"cb"),
   347 => (x"9d",x"4d",x"70",x"86"),
   348 => (x"87",x"c3",x"c3",x"02"),
   349 => (x"bf",x"c2",x"ed",x"c2"),
   350 => (x"fe",x"49",x"6e",x"4c"),
   351 => (x"ff",x"87",x"f7",x"df"),
   352 => (x"c5",x"c8",x"48",x"d0"),
   353 => (x"7b",x"d6",x"c1",x"78"),
   354 => (x"7b",x"15",x"4a",x"c0"),
   355 => (x"e0",x"c0",x"82",x"c1"),
   356 => (x"f5",x"04",x"aa",x"b7"),
   357 => (x"48",x"d0",x"ff",x"87"),
   358 => (x"c5",x"c8",x"78",x"c4"),
   359 => (x"7b",x"d3",x"c1",x"78"),
   360 => (x"78",x"c4",x"7b",x"c1"),
   361 => (x"c1",x"02",x"9c",x"74"),
   362 => (x"db",x"c2",x"87",x"fc"),
   363 => (x"c0",x"c8",x"7e",x"d6"),
   364 => (x"b7",x"c0",x"8c",x"4d"),
   365 => (x"87",x"c6",x"03",x"ac"),
   366 => (x"4d",x"a4",x"c0",x"c8"),
   367 => (x"e8",x"c2",x"4c",x"c0"),
   368 => (x"49",x"bf",x"97",x"c7"),
   369 => (x"d2",x"02",x"99",x"d0"),
   370 => (x"c2",x"1e",x"c0",x"87"),
   371 => (x"fe",x"49",x"fa",x"ec"),
   372 => (x"c4",x"87",x"cc",x"cd"),
   373 => (x"4a",x"49",x"70",x"86"),
   374 => (x"c2",x"87",x"ef",x"c0"),
   375 => (x"c2",x"1e",x"d6",x"db"),
   376 => (x"fe",x"49",x"fa",x"ec"),
   377 => (x"c4",x"87",x"f8",x"cc"),
   378 => (x"4a",x"49",x"70",x"86"),
   379 => (x"c8",x"48",x"d0",x"ff"),
   380 => (x"d4",x"c1",x"78",x"c5"),
   381 => (x"bf",x"97",x"6e",x"7b"),
   382 => (x"c1",x"48",x"6e",x"7b"),
   383 => (x"c1",x"7e",x"70",x"80"),
   384 => (x"f0",x"ff",x"05",x"8d"),
   385 => (x"48",x"d0",x"ff",x"87"),
   386 => (x"9a",x"72",x"78",x"c4"),
   387 => (x"c0",x"87",x"c5",x"05"),
   388 => (x"87",x"e5",x"c0",x"48"),
   389 => (x"ec",x"c2",x"1e",x"c1"),
   390 => (x"ca",x"fe",x"49",x"fa"),
   391 => (x"86",x"c4",x"87",x"e0"),
   392 => (x"fe",x"05",x"9c",x"74"),
   393 => (x"d0",x"ff",x"87",x"c4"),
   394 => (x"78",x"c5",x"c8",x"48"),
   395 => (x"c0",x"7b",x"d3",x"c1"),
   396 => (x"c1",x"78",x"c4",x"7b"),
   397 => (x"c0",x"87",x"c2",x"48"),
   398 => (x"4d",x"26",x"26",x"48"),
   399 => (x"4b",x"26",x"4c",x"26"),
   400 => (x"5e",x"0e",x"4f",x"26"),
   401 => (x"71",x"0e",x"5c",x"5b"),
   402 => (x"02",x"66",x"cc",x"4b"),
   403 => (x"c0",x"4c",x"87",x"d8"),
   404 => (x"d8",x"02",x"8c",x"f0"),
   405 => (x"c1",x"4a",x"74",x"87"),
   406 => (x"87",x"d1",x"02",x"8a"),
   407 => (x"87",x"cd",x"02",x"8a"),
   408 => (x"87",x"c9",x"02",x"8a"),
   409 => (x"49",x"73",x"87",x"d7"),
   410 => (x"d0",x"87",x"ea",x"fb"),
   411 => (x"c0",x"1e",x"74",x"87"),
   412 => (x"87",x"e0",x"f9",x"49"),
   413 => (x"49",x"73",x"1e",x"74"),
   414 => (x"c8",x"87",x"d9",x"f9"),
   415 => (x"87",x"fc",x"fe",x"86"),
   416 => (x"da",x"c2",x"1e",x"00"),
   417 => (x"c1",x"49",x"bf",x"ea"),
   418 => (x"ee",x"da",x"c2",x"b9"),
   419 => (x"48",x"d4",x"ff",x"59"),
   420 => (x"ff",x"78",x"ff",x"c3"),
   421 => (x"e1",x"c8",x"48",x"d0"),
   422 => (x"48",x"d4",x"ff",x"78"),
   423 => (x"31",x"c4",x"78",x"c1"),
   424 => (x"d0",x"ff",x"78",x"71"),
   425 => (x"78",x"e0",x"c0",x"48"),
   426 => (x"00",x"00",x"4f",x"26"),
   427 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

