library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d0edc287",
    12 => x"86c0c64e",
    13 => x"49d0edc2",
    14 => x"48f0dac2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087dbdb",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"66c41e4f",
    50 => x"ff48114a",
    51 => x"c17808d4",
    52 => x"87f5058a",
    53 => x"c41e4f26",
    54 => x"d4ff4a66",
    55 => x"78ffc348",
    56 => x"8ac15168",
    57 => x"2687f305",
    58 => x"1e731e4f",
    59 => x"c34bd4ff",
    60 => x"4a6b7bff",
    61 => x"6b7bffc3",
    62 => x"7232c849",
    63 => x"7bffc3b1",
    64 => x"31c84a6b",
    65 => x"ffc3b271",
    66 => x"c8496b7b",
    67 => x"71b17232",
    68 => x"2687c448",
    69 => x"264c264d",
    70 => x"0e4f264b",
    71 => x"5d5c5b5e",
    72 => x"ff4a710e",
    73 => x"49724cd4",
    74 => x"7199ffc3",
    75 => x"f0dac27c",
    76 => x"87c805bf",
    77 => x"c94866d0",
    78 => x"58a6d430",
    79 => x"d84966d0",
    80 => x"99ffc329",
    81 => x"66d07c71",
    82 => x"c329d049",
    83 => x"7c7199ff",
    84 => x"c84966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"99ffc349",
    88 => x"49727c71",
    89 => x"ffc329d0",
    90 => x"6c7c7199",
    91 => x"fff0c94b",
    92 => x"abffc34d",
    93 => x"c387d005",
    94 => x"4b6c7cff",
    95 => x"c6028dc1",
    96 => x"abffc387",
    97 => x"7387f002",
    98 => x"87c7fe48",
    99 => x"ff49c01e",
   100 => x"ffc348d4",
   101 => x"c381c178",
   102 => x"04a9b7c8",
   103 => x"4f2687f1",
   104 => x"e71e731e",
   105 => x"dff8c487",
   106 => x"c01ec04b",
   107 => x"f7c1f0ff",
   108 => x"87e7fd49",
   109 => x"a8c186c4",
   110 => x"87eac005",
   111 => x"c348d4ff",
   112 => x"c0c178ff",
   113 => x"c0c0c0c0",
   114 => x"f0e1c01e",
   115 => x"fd49e9c1",
   116 => x"86c487c9",
   117 => x"ca059870",
   118 => x"48d4ff87",
   119 => x"c178ffc3",
   120 => x"fe87cb48",
   121 => x"8bc187e6",
   122 => x"87fdfe05",
   123 => x"e6fc48c0",
   124 => x"1e731e87",
   125 => x"c348d4ff",
   126 => x"4bd378ff",
   127 => x"ffc01ec0",
   128 => x"49c1c1f0",
   129 => x"c487d4fc",
   130 => x"05987086",
   131 => x"d4ff87ca",
   132 => x"78ffc348",
   133 => x"87cb48c1",
   134 => x"c187f1fd",
   135 => x"dbff058b",
   136 => x"fb48c087",
   137 => x"5e0e87f1",
   138 => x"ff0e5c5b",
   139 => x"dbfd4cd4",
   140 => x"1eeac687",
   141 => x"c1f0e1c0",
   142 => x"defb49c8",
   143 => x"c186c487",
   144 => x"87c802a8",
   145 => x"c087eafe",
   146 => x"87e2c148",
   147 => x"7087dafa",
   148 => x"ffffcf49",
   149 => x"a9eac699",
   150 => x"fe87c802",
   151 => x"48c087d3",
   152 => x"c387cbc1",
   153 => x"f1c07cff",
   154 => x"87f4fc4b",
   155 => x"c0029870",
   156 => x"1ec087eb",
   157 => x"c1f0ffc0",
   158 => x"defa49fa",
   159 => x"7086c487",
   160 => x"87d90598",
   161 => x"6c7cffc3",
   162 => x"7cffc349",
   163 => x"c17c7c7c",
   164 => x"c40299c0",
   165 => x"d548c187",
   166 => x"d148c087",
   167 => x"05abc287",
   168 => x"48c087c4",
   169 => x"8bc187c8",
   170 => x"87fdfe05",
   171 => x"e4f948c0",
   172 => x"1e731e87",
   173 => x"48f0dac2",
   174 => x"4bc778c1",
   175 => x"c248d0ff",
   176 => x"87c8fb78",
   177 => x"c348d0ff",
   178 => x"c01ec078",
   179 => x"c0c1d0e5",
   180 => x"87c7f949",
   181 => x"a8c186c4",
   182 => x"4b87c105",
   183 => x"c505abc2",
   184 => x"c048c087",
   185 => x"8bc187f9",
   186 => x"87d0ff05",
   187 => x"c287f7fc",
   188 => x"7058f4da",
   189 => x"87cd0598",
   190 => x"ffc01ec1",
   191 => x"49d0c1f0",
   192 => x"c487d8f8",
   193 => x"48d4ff86",
   194 => x"c478ffc3",
   195 => x"dac287e0",
   196 => x"d0ff58f8",
   197 => x"ff78c248",
   198 => x"ffc348d4",
   199 => x"f748c178",
   200 => x"5e0e87f5",
   201 => x"0e5d5c5b",
   202 => x"ffc34a71",
   203 => x"4cd4ff4d",
   204 => x"d0ff7c75",
   205 => x"78c3c448",
   206 => x"1e727c75",
   207 => x"c1f0ffc0",
   208 => x"d6f749d8",
   209 => x"7086c487",
   210 => x"87c50298",
   211 => x"f0c048c0",
   212 => x"c37c7587",
   213 => x"c0c87cfe",
   214 => x"4966d41e",
   215 => x"c487e6f5",
   216 => x"757c7586",
   217 => x"d87c757c",
   218 => x"754be0da",
   219 => x"99496c7c",
   220 => x"c187c505",
   221 => x"87f3058b",
   222 => x"d0ff7c75",
   223 => x"c178c248",
   224 => x"87cff648",
   225 => x"4ad4ff1e",
   226 => x"c448d0ff",
   227 => x"ffc378d1",
   228 => x"0589c17a",
   229 => x"4f2687f8",
   230 => x"711e731e",
   231 => x"cdeec54b",
   232 => x"d4ff4adf",
   233 => x"78ffc348",
   234 => x"fec34868",
   235 => x"87c502a8",
   236 => x"ed058ac1",
   237 => x"059a7287",
   238 => x"48c087c5",
   239 => x"7387eac0",
   240 => x"87cc029b",
   241 => x"731e66c8",
   242 => x"87caf449",
   243 => x"87c686c4",
   244 => x"fe4966c8",
   245 => x"d4ff87ee",
   246 => x"78ffc348",
   247 => x"059b7378",
   248 => x"d0ff87c5",
   249 => x"c178d048",
   250 => x"87ebf448",
   251 => x"711e731e",
   252 => x"ff4bc04a",
   253 => x"ffc348d4",
   254 => x"48d0ff78",
   255 => x"ff78c3c4",
   256 => x"ffc348d4",
   257 => x"c01e7278",
   258 => x"d1c1f0ff",
   259 => x"87cbf449",
   260 => x"987086c4",
   261 => x"c887cd05",
   262 => x"66cc1ec0",
   263 => x"87f8fd49",
   264 => x"4b7086c4",
   265 => x"c248d0ff",
   266 => x"f3487378",
   267 => x"5e0e87e9",
   268 => x"0e5d5c5b",
   269 => x"ffc01ec0",
   270 => x"49c9c1f0",
   271 => x"d287dcf3",
   272 => x"f8dac21e",
   273 => x"87d0fd49",
   274 => x"4cc086c8",
   275 => x"b7d284c1",
   276 => x"87f804ac",
   277 => x"97f8dac2",
   278 => x"c0c349bf",
   279 => x"a9c0c199",
   280 => x"87e7c005",
   281 => x"97ffdac2",
   282 => x"31d049bf",
   283 => x"97c0dbc2",
   284 => x"32c84abf",
   285 => x"dbc2b172",
   286 => x"4abf97c1",
   287 => x"cf4c71b1",
   288 => x"9cffffff",
   289 => x"34ca84c1",
   290 => x"c287e7c1",
   291 => x"bf97c1db",
   292 => x"c631c149",
   293 => x"c2dbc299",
   294 => x"c74abf97",
   295 => x"b1722ab7",
   296 => x"97fddac2",
   297 => x"cf4d4abf",
   298 => x"fedac29d",
   299 => x"c34abf97",
   300 => x"c232ca9a",
   301 => x"bf97ffda",
   302 => x"7333c24b",
   303 => x"c0dbc2b2",
   304 => x"c34bbf97",
   305 => x"b7c69bc0",
   306 => x"c2b2732b",
   307 => x"7148c181",
   308 => x"c1497030",
   309 => x"70307548",
   310 => x"c14c724d",
   311 => x"c8947184",
   312 => x"06adb7c0",
   313 => x"34c187cc",
   314 => x"c0c82db7",
   315 => x"ff01adb7",
   316 => x"487487f4",
   317 => x"0e87dcf0",
   318 => x"5d5c5b5e",
   319 => x"c286f80e",
   320 => x"c048dee3",
   321 => x"d6dbc278",
   322 => x"fb49c01e",
   323 => x"86c487de",
   324 => x"c5059870",
   325 => x"c948c087",
   326 => x"4dc087ce",
   327 => x"f2c07ec1",
   328 => x"c249bfc1",
   329 => x"714accdc",
   330 => x"fdec4bc8",
   331 => x"05987087",
   332 => x"7ec087c2",
   333 => x"bffdf1c0",
   334 => x"e8dcc249",
   335 => x"4bc8714a",
   336 => x"7087e7ec",
   337 => x"87c20598",
   338 => x"026e7ec0",
   339 => x"c287fdc0",
   340 => x"4dbfdce2",
   341 => x"9fd4e3c2",
   342 => x"c5487ebf",
   343 => x"05a8ead6",
   344 => x"e2c287c7",
   345 => x"ce4dbfdc",
   346 => x"ca486e87",
   347 => x"02a8d5e9",
   348 => x"48c087c5",
   349 => x"c287f1c7",
   350 => x"751ed6db",
   351 => x"87ecf949",
   352 => x"987086c4",
   353 => x"c087c505",
   354 => x"87dcc748",
   355 => x"bffdf1c0",
   356 => x"e8dcc249",
   357 => x"4bc8714a",
   358 => x"7087cfeb",
   359 => x"87c80598",
   360 => x"48dee3c2",
   361 => x"87da78c1",
   362 => x"bfc1f2c0",
   363 => x"ccdcc249",
   364 => x"4bc8714a",
   365 => x"7087f3ea",
   366 => x"c5c00298",
   367 => x"c648c087",
   368 => x"e3c287e6",
   369 => x"49bf97d4",
   370 => x"05a9d5c1",
   371 => x"c287cdc0",
   372 => x"bf97d5e3",
   373 => x"a9eac249",
   374 => x"87c5c002",
   375 => x"c7c648c0",
   376 => x"d6dbc287",
   377 => x"487ebf97",
   378 => x"02a8e9c3",
   379 => x"6e87cec0",
   380 => x"a8ebc348",
   381 => x"87c5c002",
   382 => x"ebc548c0",
   383 => x"e1dbc287",
   384 => x"9949bf97",
   385 => x"87ccc005",
   386 => x"97e2dbc2",
   387 => x"a9c249bf",
   388 => x"87c5c002",
   389 => x"cfc548c0",
   390 => x"e3dbc287",
   391 => x"c248bf97",
   392 => x"7058dae3",
   393 => x"88c1484c",
   394 => x"58dee3c2",
   395 => x"97e4dbc2",
   396 => x"817549bf",
   397 => x"97e5dbc2",
   398 => x"32c84abf",
   399 => x"c27ea172",
   400 => x"6e48ebe7",
   401 => x"e6dbc278",
   402 => x"c848bf97",
   403 => x"e3c258a6",
   404 => x"c202bfde",
   405 => x"f1c087d4",
   406 => x"c249bffd",
   407 => x"714ae8dc",
   408 => x"c5e84bc8",
   409 => x"02987087",
   410 => x"c087c5c0",
   411 => x"87f8c348",
   412 => x"bfd6e3c2",
   413 => x"ffe7c24c",
   414 => x"fbdbc25c",
   415 => x"c849bf97",
   416 => x"fadbc231",
   417 => x"a14abf97",
   418 => x"fcdbc249",
   419 => x"d04abf97",
   420 => x"49a17232",
   421 => x"97fddbc2",
   422 => x"32d84abf",
   423 => x"c449a172",
   424 => x"e7c29166",
   425 => x"c281bfeb",
   426 => x"c259f3e7",
   427 => x"bf97c3dc",
   428 => x"c232c84a",
   429 => x"bf97c2dc",
   430 => x"c24aa24b",
   431 => x"bf97c4dc",
   432 => x"7333d04b",
   433 => x"dcc24aa2",
   434 => x"4bbf97c5",
   435 => x"33d89bcf",
   436 => x"c24aa273",
   437 => x"c25af7e7",
   438 => x"4abff3e7",
   439 => x"92748ac2",
   440 => x"48f7e7c2",
   441 => x"c178a172",
   442 => x"dbc287ca",
   443 => x"49bf97e8",
   444 => x"dbc231c8",
   445 => x"4abf97e7",
   446 => x"e3c249a1",
   447 => x"e3c259e6",
   448 => x"c549bfe2",
   449 => x"81ffc731",
   450 => x"e7c229c9",
   451 => x"dbc259ff",
   452 => x"4abf97ed",
   453 => x"dbc232c8",
   454 => x"4bbf97ec",
   455 => x"66c44aa2",
   456 => x"c2826e92",
   457 => x"c25afbe7",
   458 => x"c048f3e7",
   459 => x"efe7c278",
   460 => x"78a17248",
   461 => x"48ffe7c2",
   462 => x"bff3e7c2",
   463 => x"c3e8c278",
   464 => x"f7e7c248",
   465 => x"e3c278bf",
   466 => x"c002bfde",
   467 => x"487487c9",
   468 => x"7e7030c4",
   469 => x"c287c9c0",
   470 => x"48bffbe7",
   471 => x"7e7030c4",
   472 => x"48e2e3c2",
   473 => x"48c1786e",
   474 => x"4d268ef8",
   475 => x"4b264c26",
   476 => x"5e0e4f26",
   477 => x"0e5d5c5b",
   478 => x"e3c24a71",
   479 => x"cb02bfde",
   480 => x"c74b7287",
   481 => x"c14c722b",
   482 => x"87c99cff",
   483 => x"2bc84b72",
   484 => x"ffc34c72",
   485 => x"ebe7c29c",
   486 => x"f1c083bf",
   487 => x"02abbff9",
   488 => x"f1c087d9",
   489 => x"dbc25bfd",
   490 => x"49731ed6",
   491 => x"c487fdf0",
   492 => x"05987086",
   493 => x"48c087c5",
   494 => x"c287e6c0",
   495 => x"02bfdee3",
   496 => x"497487d2",
   497 => x"dbc291c4",
   498 => x"4d6981d6",
   499 => x"ffffffcf",
   500 => x"87cb9dff",
   501 => x"91c24974",
   502 => x"81d6dbc2",
   503 => x"754d699f",
   504 => x"87c6fe48",
   505 => x"5c5b5e0e",
   506 => x"711e0e5d",
   507 => x"c11ec04d",
   508 => x"87eeca49",
   509 => x"4c7086c4",
   510 => x"c0c1029c",
   511 => x"e6e3c287",
   512 => x"e149754a",
   513 => x"987087c9",
   514 => x"87f1c002",
   515 => x"49754a74",
   516 => x"efe14bcb",
   517 => x"02987087",
   518 => x"c087e2c0",
   519 => x"029c741e",
   520 => x"a6c487c7",
   521 => x"c578c048",
   522 => x"48a6c487",
   523 => x"66c478c1",
   524 => x"87eec949",
   525 => x"4c7086c4",
   526 => x"c0ff059c",
   527 => x"26487487",
   528 => x"0e87e7fc",
   529 => x"5d5c5b5e",
   530 => x"4b711e0e",
   531 => x"87c5059b",
   532 => x"e5c148c0",
   533 => x"4da3c887",
   534 => x"66d47dc0",
   535 => x"d487c702",
   536 => x"05bf9766",
   537 => x"48c087c5",
   538 => x"d487cfc1",
   539 => x"f3fd4966",
   540 => x"9c4c7087",
   541 => x"87c0c102",
   542 => x"6949a4dc",
   543 => x"49a4da7d",
   544 => x"9f4aa3c4",
   545 => x"e3c27a69",
   546 => x"d202bfde",
   547 => x"49a4d487",
   548 => x"c049699f",
   549 => x"7199ffff",
   550 => x"7030d048",
   551 => x"c087c27e",
   552 => x"48496e7e",
   553 => x"7a70806a",
   554 => x"a3cc7bc0",
   555 => x"d0796a49",
   556 => x"79c049a3",
   557 => x"87c24874",
   558 => x"fa2648c0",
   559 => x"5e0e87ec",
   560 => x"0e5d5c5b",
   561 => x"f1c04c71",
   562 => x"78ff48f9",
   563 => x"c1029c74",
   564 => x"a4c887ca",
   565 => x"c1026949",
   566 => x"66d087c2",
   567 => x"82496c4a",
   568 => x"d05aa6d4",
   569 => x"c2b94d66",
   570 => x"4abfdae3",
   571 => x"9972baff",
   572 => x"c0029971",
   573 => x"a4c487e4",
   574 => x"f9496b4b",
   575 => x"7b7087f4",
   576 => x"bfd6e3c2",
   577 => x"71816c49",
   578 => x"c2b9757c",
   579 => x"4abfdae3",
   580 => x"9972baff",
   581 => x"ff059971",
   582 => x"7c7587dc",
   583 => x"1e87cbf9",
   584 => x"4b711e73",
   585 => x"87c7029b",
   586 => x"6949a3c8",
   587 => x"c087c505",
   588 => x"87ebc048",
   589 => x"bfefe7c2",
   590 => x"49a3c44a",
   591 => x"89c24969",
   592 => x"bfd6e3c2",
   593 => x"4aa27191",
   594 => x"bfdae3c2",
   595 => x"71996b49",
   596 => x"66c84aa2",
   597 => x"ea49721e",
   598 => x"86c487d2",
   599 => x"f8484970",
   600 => x"731e87cc",
   601 => x"9b4b711e",
   602 => x"c887c702",
   603 => x"056949a3",
   604 => x"48c087c5",
   605 => x"c287ebc0",
   606 => x"4abfefe7",
   607 => x"6949a3c4",
   608 => x"c289c249",
   609 => x"91bfd6e3",
   610 => x"c24aa271",
   611 => x"49bfdae3",
   612 => x"a271996b",
   613 => x"1e66c84a",
   614 => x"c5e64972",
   615 => x"7086c487",
   616 => x"c9f74849",
   617 => x"5b5e0e87",
   618 => x"1e0e5d5c",
   619 => x"66d44b71",
   620 => x"732cc94c",
   621 => x"cfc1029b",
   622 => x"49a3c887",
   623 => x"c7c10269",
   624 => x"4da3d087",
   625 => x"c27d66d4",
   626 => x"49bfdae3",
   627 => x"4a6bb9ff",
   628 => x"ac717e99",
   629 => x"c087cd03",
   630 => x"a3cc7d7b",
   631 => x"49a3c44a",
   632 => x"87c2796a",
   633 => x"9c748c72",
   634 => x"4987dd02",
   635 => x"fb49731e",
   636 => x"86c487cc",
   637 => x"c74966d4",
   638 => x"cb0299ff",
   639 => x"d6dbc287",
   640 => x"fc49731e",
   641 => x"86c487d9",
   642 => x"87def526",
   643 => x"711e731e",
   644 => x"c0029b4b",
   645 => x"e8c287e4",
   646 => x"4a735bc3",
   647 => x"e3c28ac2",
   648 => x"9249bfd6",
   649 => x"bfefe7c2",
   650 => x"c2807248",
   651 => x"7158c7e8",
   652 => x"c230c448",
   653 => x"c058e6e3",
   654 => x"e7c287ed",
   655 => x"e7c248ff",
   656 => x"c278bff3",
   657 => x"c248c3e8",
   658 => x"78bff7e7",
   659 => x"bfdee3c2",
   660 => x"c287c902",
   661 => x"49bfd6e3",
   662 => x"87c731c4",
   663 => x"bffbe7c2",
   664 => x"c231c449",
   665 => x"f459e6e3",
   666 => x"5e0e87c4",
   667 => x"710e5c5b",
   668 => x"724bc04a",
   669 => x"e1c0029a",
   670 => x"49a2da87",
   671 => x"c24b699f",
   672 => x"02bfdee3",
   673 => x"a2d487cf",
   674 => x"49699f49",
   675 => x"ffffc04c",
   676 => x"c234d09c",
   677 => x"744cc087",
   678 => x"4973b349",
   679 => x"f387edfd",
   680 => x"5e0e87ca",
   681 => x"0e5d5c5b",
   682 => x"4a7186f4",
   683 => x"9a727ec0",
   684 => x"c287d802",
   685 => x"c048d2db",
   686 => x"cadbc278",
   687 => x"c3e8c248",
   688 => x"dbc278bf",
   689 => x"e7c248ce",
   690 => x"c278bfff",
   691 => x"c048f3e3",
   692 => x"e2e3c250",
   693 => x"dbc249bf",
   694 => x"714abfd2",
   695 => x"ffc303aa",
   696 => x"cf497287",
   697 => x"e0c00599",
   698 => x"d6dbc287",
   699 => x"cadbc21e",
   700 => x"dbc249bf",
   701 => x"a1c148ca",
   702 => x"efe37178",
   703 => x"c086c487",
   704 => x"c248f5f1",
   705 => x"cc78d6db",
   706 => x"f5f1c087",
   707 => x"e0c048bf",
   708 => x"f9f1c080",
   709 => x"d2dbc258",
   710 => x"80c148bf",
   711 => x"58d6dbc2",
   712 => x"000c7527",
   713 => x"bf97bf00",
   714 => x"c2029d4d",
   715 => x"e5c387e2",
   716 => x"dbc202ad",
   717 => x"f5f1c087",
   718 => x"a3cb4bbf",
   719 => x"cf4c1149",
   720 => x"d2c105ac",
   721 => x"df497587",
   722 => x"cd89c199",
   723 => x"e6e3c291",
   724 => x"4aa3c181",
   725 => x"a3c35112",
   726 => x"c551124a",
   727 => x"51124aa3",
   728 => x"124aa3c7",
   729 => x"4aa3c951",
   730 => x"a3ce5112",
   731 => x"d051124a",
   732 => x"51124aa3",
   733 => x"124aa3d2",
   734 => x"4aa3d451",
   735 => x"a3d65112",
   736 => x"d851124a",
   737 => x"51124aa3",
   738 => x"124aa3dc",
   739 => x"4aa3de51",
   740 => x"7ec15112",
   741 => x"7487f9c0",
   742 => x"0599c849",
   743 => x"7487eac0",
   744 => x"0599d049",
   745 => x"66dc87d0",
   746 => x"87cac002",
   747 => x"66dc4973",
   748 => x"0298700f",
   749 => x"056e87d3",
   750 => x"c287c6c0",
   751 => x"c048e6e3",
   752 => x"f5f1c050",
   753 => x"e7c248bf",
   754 => x"f3e3c287",
   755 => x"7e50c048",
   756 => x"bfe2e3c2",
   757 => x"d2dbc249",
   758 => x"aa714abf",
   759 => x"87c1fc04",
   760 => x"bfc3e8c2",
   761 => x"87c8c005",
   762 => x"bfdee3c2",
   763 => x"87fec102",
   764 => x"48f9f1c0",
   765 => x"dbc278ff",
   766 => x"ed49bfce",
   767 => x"497087f4",
   768 => x"59d2dbc2",
   769 => x"c248a6c4",
   770 => x"78bfcedb",
   771 => x"bfdee3c2",
   772 => x"87d8c002",
   773 => x"cf4966c4",
   774 => x"f8ffffff",
   775 => x"c002a999",
   776 => x"4dc087c5",
   777 => x"c187e1c0",
   778 => x"87dcc04d",
   779 => x"cf4966c4",
   780 => x"a999f8ff",
   781 => x"87c8c002",
   782 => x"c048a6c8",
   783 => x"87c5c078",
   784 => x"c148a6c8",
   785 => x"4d66c878",
   786 => x"c0059d75",
   787 => x"66c487e0",
   788 => x"c289c249",
   789 => x"4abfd6e3",
   790 => x"efe7c291",
   791 => x"dbc24abf",
   792 => x"a17248ca",
   793 => x"d2dbc278",
   794 => x"f978c048",
   795 => x"48c087e3",
   796 => x"f5eb8ef4",
   797 => x"00000087",
   798 => x"ffffff00",
   799 => x"000c85ff",
   800 => x"000c8e00",
   801 => x"54414600",
   802 => x"20203233",
   803 => x"41460020",
   804 => x"20363154",
   805 => x"1e002020",
   806 => x"c348d4ff",
   807 => x"486878ff",
   808 => x"ff1e4f26",
   809 => x"ffc348d4",
   810 => x"48d0ff78",
   811 => x"ff78e1c8",
   812 => x"78d448d4",
   813 => x"48c7e8c2",
   814 => x"50bfd4ff",
   815 => x"ff1e4f26",
   816 => x"e0c048d0",
   817 => x"1e4f2678",
   818 => x"7087ccff",
   819 => x"c6029949",
   820 => x"a9fbc087",
   821 => x"7187f105",
   822 => x"0e4f2648",
   823 => x"0e5c5b5e",
   824 => x"4cc04b71",
   825 => x"7087f0fe",
   826 => x"c0029949",
   827 => x"ecc087f9",
   828 => x"f2c002a9",
   829 => x"a9fbc087",
   830 => x"87ebc002",
   831 => x"acb766cc",
   832 => x"d087c703",
   833 => x"87c20266",
   834 => x"99715371",
   835 => x"c187c202",
   836 => x"87c3fe84",
   837 => x"02994970",
   838 => x"ecc087cd",
   839 => x"87c702a9",
   840 => x"05a9fbc0",
   841 => x"d087d5ff",
   842 => x"87c30266",
   843 => x"c07b97c0",
   844 => x"c405a9ec",
   845 => x"c54a7487",
   846 => x"c04a7487",
   847 => x"48728a0a",
   848 => x"4d2687c2",
   849 => x"4b264c26",
   850 => x"fd1e4f26",
   851 => x"497087c9",
   852 => x"a9b7f0c0",
   853 => x"c087ca04",
   854 => x"01a9b7f9",
   855 => x"f0c087c3",
   856 => x"b7c1c189",
   857 => x"87ca04a9",
   858 => x"a9b7dac1",
   859 => x"c087c301",
   860 => x"487189f7",
   861 => x"5e0e4f26",
   862 => x"710e5c5b",
   863 => x"4cd4ff4a",
   864 => x"eac04972",
   865 => x"9b4b7087",
   866 => x"c187c202",
   867 => x"48d0ff8b",
   868 => x"c178c5c8",
   869 => x"49737cd5",
   870 => x"dac231c6",
   871 => x"4abf97c0",
   872 => x"70b07148",
   873 => x"48d0ff7c",
   874 => x"487378c4",
   875 => x"0e87d5fe",
   876 => x"5d5c5b5e",
   877 => x"7186f80e",
   878 => x"fb7ec04c",
   879 => x"4bc087e4",
   880 => x"97dcf9c0",
   881 => x"a9c049bf",
   882 => x"fb87cf04",
   883 => x"83c187f9",
   884 => x"97dcf9c0",
   885 => x"06ab49bf",
   886 => x"f9c087f1",
   887 => x"02bf97dc",
   888 => x"f2fa87cf",
   889 => x"99497087",
   890 => x"c087c602",
   891 => x"f105a9ec",
   892 => x"fa4bc087",
   893 => x"4d7087e1",
   894 => x"c887dcfa",
   895 => x"d6fa58a6",
   896 => x"c14a7087",
   897 => x"49a4c883",
   898 => x"ad496997",
   899 => x"c087c702",
   900 => x"c005adff",
   901 => x"a4c987e7",
   902 => x"49699749",
   903 => x"02a966c4",
   904 => x"c04887c7",
   905 => x"d405a8ff",
   906 => x"49a4ca87",
   907 => x"aa496997",
   908 => x"c087c602",
   909 => x"c405aaff",
   910 => x"d07ec187",
   911 => x"adecc087",
   912 => x"c087c602",
   913 => x"c405adfb",
   914 => x"c14bc087",
   915 => x"fe026e7e",
   916 => x"e9f987e1",
   917 => x"f8487387",
   918 => x"87e6fb8e",
   919 => x"5b5e0e00",
   920 => x"1e0e5d5c",
   921 => x"4cc04b71",
   922 => x"c004ab4d",
   923 => x"f6c087e8",
   924 => x"9d751eef",
   925 => x"c087c402",
   926 => x"c187c24a",
   927 => x"f049724a",
   928 => x"86c487e0",
   929 => x"84c17e70",
   930 => x"87c2056e",
   931 => x"85c14c73",
   932 => x"ff06ac73",
   933 => x"486e87d8",
   934 => x"264d2626",
   935 => x"264b264c",
   936 => x"5b5e0e4f",
   937 => x"1e0e5d5c",
   938 => x"de494c71",
   939 => x"e1e8c291",
   940 => x"9785714d",
   941 => x"ddc1026d",
   942 => x"cce8c287",
   943 => x"82744abf",
   944 => x"d8fe4972",
   945 => x"6e7e7087",
   946 => x"87f3c002",
   947 => x"4bd4e8c2",
   948 => x"49cb4a6e",
   949 => x"87d0c7ff",
   950 => x"93cb4b74",
   951 => x"83caddc1",
   952 => x"fcc083c4",
   953 => x"49747bda",
   954 => x"87ebc2c1",
   955 => x"e8c27b75",
   956 => x"49bf97e0",
   957 => x"d4e8c21e",
   958 => x"c5ddc149",
   959 => x"7486c487",
   960 => x"d2c2c149",
   961 => x"c149c087",
   962 => x"c287f1c3",
   963 => x"c048c8e8",
   964 => x"dd49c178",
   965 => x"fd2687cb",
   966 => x"6f4c87ff",
   967 => x"6e696461",
   968 => x"2e2e2e67",
   969 => x"5b5e0e00",
   970 => x"4b710e5c",
   971 => x"cce8c24a",
   972 => x"497282bf",
   973 => x"7087e6fc",
   974 => x"c4029c4c",
   975 => x"e9ec4987",
   976 => x"cce8c287",
   977 => x"c178c048",
   978 => x"87d5dc49",
   979 => x"0e87ccfd",
   980 => x"5d5c5b5e",
   981 => x"c286f40e",
   982 => x"c04dd6db",
   983 => x"48a6c44c",
   984 => x"e8c278c0",
   985 => x"c049bfcc",
   986 => x"c1c106a9",
   987 => x"d6dbc287",
   988 => x"c0029848",
   989 => x"f6c087f8",
   990 => x"66c81eef",
   991 => x"c487c702",
   992 => x"78c048a6",
   993 => x"a6c487c5",
   994 => x"c478c148",
   995 => x"d1ec4966",
   996 => x"7086c487",
   997 => x"c484c14d",
   998 => x"80c14866",
   999 => x"c258a6c8",
  1000 => x"49bfcce8",
  1001 => x"87c603ac",
  1002 => x"ff059d75",
  1003 => x"4cc087c8",
  1004 => x"c3029d75",
  1005 => x"f6c087e0",
  1006 => x"66c81eef",
  1007 => x"cc87c702",
  1008 => x"78c048a6",
  1009 => x"a6cc87c5",
  1010 => x"cc78c148",
  1011 => x"d1eb4966",
  1012 => x"7086c487",
  1013 => x"c2026e7e",
  1014 => x"496e87e9",
  1015 => x"699781cb",
  1016 => x"0299d049",
  1017 => x"c087d6c1",
  1018 => x"744ae5fc",
  1019 => x"c191cb49",
  1020 => x"7281cadd",
  1021 => x"c381c879",
  1022 => x"497451ff",
  1023 => x"e8c291de",
  1024 => x"85714de1",
  1025 => x"7d97c1c2",
  1026 => x"c049a5c1",
  1027 => x"e3c251e0",
  1028 => x"02bf97e6",
  1029 => x"84c187d2",
  1030 => x"c24ba5c2",
  1031 => x"db4ae6e3",
  1032 => x"c3c2ff49",
  1033 => x"87dbc187",
  1034 => x"c049a5cd",
  1035 => x"c284c151",
  1036 => x"4a6e4ba5",
  1037 => x"c1ff49cb",
  1038 => x"c6c187ee",
  1039 => x"e1fac087",
  1040 => x"cb49744a",
  1041 => x"caddc191",
  1042 => x"c2797281",
  1043 => x"bf97e6e3",
  1044 => x"7487d802",
  1045 => x"c191de49",
  1046 => x"e1e8c284",
  1047 => x"c283714b",
  1048 => x"dd4ae6e3",
  1049 => x"ffc0ff49",
  1050 => x"7487d887",
  1051 => x"c293de4b",
  1052 => x"cb83e1e8",
  1053 => x"51c049a3",
  1054 => x"6e7384c1",
  1055 => x"ff49cb4a",
  1056 => x"c487e5c0",
  1057 => x"80c14866",
  1058 => x"c758a6c8",
  1059 => x"c5c003ac",
  1060 => x"fc056e87",
  1061 => x"487487e0",
  1062 => x"fcf78ef4",
  1063 => x"1e731e87",
  1064 => x"cb494b71",
  1065 => x"caddc191",
  1066 => x"4aa1c881",
  1067 => x"48c0dac2",
  1068 => x"a1c95012",
  1069 => x"dcf9c04a",
  1070 => x"ca501248",
  1071 => x"e0e8c281",
  1072 => x"c2501148",
  1073 => x"bf97e0e8",
  1074 => x"49c01e49",
  1075 => x"87f2d5c1",
  1076 => x"48c8e8c2",
  1077 => x"49c178de",
  1078 => x"2687c6d6",
  1079 => x"1e87fef6",
  1080 => x"cb494a71",
  1081 => x"caddc191",
  1082 => x"1181c881",
  1083 => x"cce8c248",
  1084 => x"cce8c258",
  1085 => x"c178c048",
  1086 => x"87e5d549",
  1087 => x"c01e4f26",
  1088 => x"f7fbc049",
  1089 => x"1e4f2687",
  1090 => x"d2029971",
  1091 => x"dfdec187",
  1092 => x"f750c048",
  1093 => x"dfc3c180",
  1094 => x"c3ddc140",
  1095 => x"c187ce78",
  1096 => x"c148dbde",
  1097 => x"fc78fcdc",
  1098 => x"fec3c180",
  1099 => x"0e4f2678",
  1100 => x"0e5c5b5e",
  1101 => x"cb4a4c71",
  1102 => x"caddc192",
  1103 => x"49a2c882",
  1104 => x"974ba2c9",
  1105 => x"971e4b6b",
  1106 => x"ca1e4969",
  1107 => x"c0491282",
  1108 => x"c087f2e6",
  1109 => x"87c9d449",
  1110 => x"f8c04974",
  1111 => x"8ef887f9",
  1112 => x"1e87f8f4",
  1113 => x"4b711e73",
  1114 => x"87c3ff49",
  1115 => x"fefe4973",
  1116 => x"87e9f487",
  1117 => x"711e731e",
  1118 => x"4aa3c64b",
  1119 => x"c187db02",
  1120 => x"87d6028a",
  1121 => x"dac1028a",
  1122 => x"c0028a87",
  1123 => x"028a87fc",
  1124 => x"8a87e1c0",
  1125 => x"c187cb02",
  1126 => x"49c787db",
  1127 => x"c187c0fd",
  1128 => x"e8c287de",
  1129 => x"c102bfcc",
  1130 => x"c14887cb",
  1131 => x"d0e8c288",
  1132 => x"87c1c158",
  1133 => x"bfd0e8c2",
  1134 => x"87f9c002",
  1135 => x"bfcce8c2",
  1136 => x"c280c148",
  1137 => x"c058d0e8",
  1138 => x"e8c287eb",
  1139 => x"c649bfcc",
  1140 => x"d0e8c289",
  1141 => x"a9b7c059",
  1142 => x"c287da03",
  1143 => x"c048cce8",
  1144 => x"c287d278",
  1145 => x"02bfd0e8",
  1146 => x"e8c287cb",
  1147 => x"c648bfcc",
  1148 => x"d0e8c280",
  1149 => x"d149c058",
  1150 => x"497387e7",
  1151 => x"87d7f6c0",
  1152 => x"0e87daf2",
  1153 => x"0e5c5b5e",
  1154 => x"66cc4c71",
  1155 => x"cb4b741e",
  1156 => x"caddc193",
  1157 => x"4aa3c483",
  1158 => x"fafe496a",
  1159 => x"c2c187da",
  1160 => x"a3c87bdd",
  1161 => x"5166d449",
  1162 => x"d849a3c9",
  1163 => x"a3ca5166",
  1164 => x"5166dc49",
  1165 => x"87e3f126",
  1166 => x"5c5b5e0e",
  1167 => x"d0ff0e5d",
  1168 => x"59a6d886",
  1169 => x"c048a6c4",
  1170 => x"c180c478",
  1171 => x"c47866c4",
  1172 => x"c478c180",
  1173 => x"c278c180",
  1174 => x"c148d0e8",
  1175 => x"c8e8c278",
  1176 => x"a8de48bf",
  1177 => x"f387cb05",
  1178 => x"497087e5",
  1179 => x"ce59a6c8",
  1180 => x"ede887f8",
  1181 => x"87cfe987",
  1182 => x"7087dce8",
  1183 => x"acfbc04c",
  1184 => x"87d0c102",
  1185 => x"c10566d4",
  1186 => x"1ec087c2",
  1187 => x"c11ec11e",
  1188 => x"c01efdde",
  1189 => x"87ebfd49",
  1190 => x"4a66d0c1",
  1191 => x"496a82c4",
  1192 => x"517481c7",
  1193 => x"1ed81ec1",
  1194 => x"81c8496a",
  1195 => x"d887ece8",
  1196 => x"66c4c186",
  1197 => x"01a8c048",
  1198 => x"a6c487c7",
  1199 => x"ce78c148",
  1200 => x"66c4c187",
  1201 => x"cc88c148",
  1202 => x"87c358a6",
  1203 => x"cc87f8e7",
  1204 => x"78c248a6",
  1205 => x"cd029c74",
  1206 => x"66c487cc",
  1207 => x"66c8c148",
  1208 => x"c1cd03a8",
  1209 => x"48a6d887",
  1210 => x"eae678c0",
  1211 => x"c14c7087",
  1212 => x"c205acd0",
  1213 => x"66d887d6",
  1214 => x"87cee97e",
  1215 => x"a6dc4970",
  1216 => x"87d3e659",
  1217 => x"ecc04c70",
  1218 => x"eac105ac",
  1219 => x"4966c487",
  1220 => x"c0c191cb",
  1221 => x"a1c48166",
  1222 => x"c84d6a4a",
  1223 => x"66d84aa1",
  1224 => x"dfc3c152",
  1225 => x"87efe579",
  1226 => x"029c4c70",
  1227 => x"fbc087d8",
  1228 => x"87d202ac",
  1229 => x"dee55574",
  1230 => x"9c4c7087",
  1231 => x"c087c702",
  1232 => x"ff05acfb",
  1233 => x"e0c087ee",
  1234 => x"55c1c255",
  1235 => x"d47d97c0",
  1236 => x"a96e4966",
  1237 => x"c487db05",
  1238 => x"66c84866",
  1239 => x"87ca04a8",
  1240 => x"c14866c4",
  1241 => x"58a6c880",
  1242 => x"66c887c8",
  1243 => x"cc88c148",
  1244 => x"e2e458a6",
  1245 => x"c14c7087",
  1246 => x"c805acd0",
  1247 => x"4866d087",
  1248 => x"a6d480c1",
  1249 => x"acd0c158",
  1250 => x"87eafd02",
  1251 => x"d448a6dc",
  1252 => x"66d87866",
  1253 => x"a866dc48",
  1254 => x"87dcc905",
  1255 => x"48a6e0c0",
  1256 => x"c478f0c0",
  1257 => x"7866cc80",
  1258 => x"78c080c4",
  1259 => x"c048747e",
  1260 => x"f0c088fb",
  1261 => x"987058a6",
  1262 => x"87d7c802",
  1263 => x"c088cb48",
  1264 => x"7058a6f0",
  1265 => x"e9c00298",
  1266 => x"88c94887",
  1267 => x"58a6f0c0",
  1268 => x"c3029870",
  1269 => x"c44887e1",
  1270 => x"a6f0c088",
  1271 => x"02987058",
  1272 => x"c14887d6",
  1273 => x"a6f0c088",
  1274 => x"02987058",
  1275 => x"c787c8c3",
  1276 => x"e0c087db",
  1277 => x"78c048a6",
  1278 => x"c14866cc",
  1279 => x"58a6d080",
  1280 => x"7087d4e2",
  1281 => x"acecc04c",
  1282 => x"c087d502",
  1283 => x"c60266e0",
  1284 => x"a6e4c087",
  1285 => x"7487c95c",
  1286 => x"88f0c048",
  1287 => x"58a6e8c0",
  1288 => x"02acecc0",
  1289 => x"eee187cc",
  1290 => x"c04c7087",
  1291 => x"ff05acec",
  1292 => x"e0c087f4",
  1293 => x"66d41e66",
  1294 => x"ecc01e49",
  1295 => x"dec11e66",
  1296 => x"66d41efd",
  1297 => x"87fbf649",
  1298 => x"1eca1ec0",
  1299 => x"cb4966dc",
  1300 => x"66d8c191",
  1301 => x"48a6d881",
  1302 => x"d878a1c4",
  1303 => x"e149bf66",
  1304 => x"86d887f9",
  1305 => x"06a8b7c0",
  1306 => x"c187c7c1",
  1307 => x"c81ede1e",
  1308 => x"e149bf66",
  1309 => x"86c887e5",
  1310 => x"c0484970",
  1311 => x"e4c08808",
  1312 => x"b7c058a6",
  1313 => x"e9c006a8",
  1314 => x"66e0c087",
  1315 => x"a8b7dd48",
  1316 => x"6e87df03",
  1317 => x"e0c049bf",
  1318 => x"e0c08166",
  1319 => x"c1496651",
  1320 => x"81bf6e81",
  1321 => x"c051c1c2",
  1322 => x"c24966e0",
  1323 => x"81bf6e81",
  1324 => x"7ec151c0",
  1325 => x"e287dcc4",
  1326 => x"e4c087d0",
  1327 => x"c9e258a6",
  1328 => x"a6e8c087",
  1329 => x"a8ecc058",
  1330 => x"87cbc005",
  1331 => x"48a6e4c0",
  1332 => x"7866e0c0",
  1333 => x"ff87c4c0",
  1334 => x"c487fcde",
  1335 => x"91cb4966",
  1336 => x"4866c0c1",
  1337 => x"7e708071",
  1338 => x"82c84a6e",
  1339 => x"81ca496e",
  1340 => x"5166e0c0",
  1341 => x"4966e4c0",
  1342 => x"e0c081c1",
  1343 => x"48c18966",
  1344 => x"49703071",
  1345 => x"977189c1",
  1346 => x"fdebc27a",
  1347 => x"e0c049bf",
  1348 => x"6a972966",
  1349 => x"9871484a",
  1350 => x"58a6f0c0",
  1351 => x"81c4496e",
  1352 => x"66dc4d69",
  1353 => x"a866d848",
  1354 => x"87c8c002",
  1355 => x"c048a6d8",
  1356 => x"87c5c078",
  1357 => x"c148a6d8",
  1358 => x"1e66d878",
  1359 => x"751ee0c0",
  1360 => x"d6deff49",
  1361 => x"7086c887",
  1362 => x"acb7c04c",
  1363 => x"87d4c106",
  1364 => x"e0c08574",
  1365 => x"75897449",
  1366 => x"ded9c14b",
  1367 => x"edfe714a",
  1368 => x"85c287c6",
  1369 => x"4866e8c0",
  1370 => x"ecc080c1",
  1371 => x"ecc058a6",
  1372 => x"81c14966",
  1373 => x"c002a970",
  1374 => x"a6d887c8",
  1375 => x"c078c048",
  1376 => x"a6d887c5",
  1377 => x"d878c148",
  1378 => x"a4c21e66",
  1379 => x"48e0c049",
  1380 => x"49708871",
  1381 => x"ff49751e",
  1382 => x"c887c0dd",
  1383 => x"a8b7c086",
  1384 => x"87c0ff01",
  1385 => x"0266e8c0",
  1386 => x"6e87d1c0",
  1387 => x"c081c949",
  1388 => x"6e5166e8",
  1389 => x"efc4c148",
  1390 => x"87ccc078",
  1391 => x"81c9496e",
  1392 => x"486e51c2",
  1393 => x"78e3c5c1",
  1394 => x"c6c07ec1",
  1395 => x"f6dbff87",
  1396 => x"6e4c7087",
  1397 => x"87f5c002",
  1398 => x"c84866c4",
  1399 => x"c004a866",
  1400 => x"66c487cb",
  1401 => x"c880c148",
  1402 => x"e0c058a6",
  1403 => x"4866c887",
  1404 => x"a6cc88c1",
  1405 => x"87d5c058",
  1406 => x"05acc6c1",
  1407 => x"cc87c8c0",
  1408 => x"80c14866",
  1409 => x"ff58a6d0",
  1410 => x"7087fcda",
  1411 => x"4866d04c",
  1412 => x"a6d480c1",
  1413 => x"029c7458",
  1414 => x"c487cbc0",
  1415 => x"c8c14866",
  1416 => x"f204a866",
  1417 => x"daff87ff",
  1418 => x"66c487d4",
  1419 => x"03a8c748",
  1420 => x"c287e5c0",
  1421 => x"c048d0e8",
  1422 => x"4966c478",
  1423 => x"c0c191cb",
  1424 => x"a1c48166",
  1425 => x"c04a6a4a",
  1426 => x"66c47952",
  1427 => x"c880c148",
  1428 => x"a8c758a6",
  1429 => x"87dbff04",
  1430 => x"e08ed0ff",
  1431 => x"203a87fb",
  1432 => x"1e731e00",
  1433 => x"029b4b71",
  1434 => x"e8c287c6",
  1435 => x"78c048cc",
  1436 => x"e8c21ec7",
  1437 => x"1e49bfcc",
  1438 => x"1ecaddc1",
  1439 => x"bfc8e8c2",
  1440 => x"87f4ee49",
  1441 => x"e8c286cc",
  1442 => x"e949bfc8",
  1443 => x"9b7387f9",
  1444 => x"c187c802",
  1445 => x"c049cadd",
  1446 => x"ff87cee5",
  1447 => x"1e87fedf",
  1448 => x"48c0dac2",
  1449 => x"dec150c0",
  1450 => x"c049bfed",
  1451 => x"c087e6fa",
  1452 => x"1e4f2648",
  1453 => x"c187e5c7",
  1454 => x"87e5fe49",
  1455 => x"87f1effe",
  1456 => x"cd029870",
  1457 => x"eef8fe87",
  1458 => x"02987087",
  1459 => x"4ac187c4",
  1460 => x"4ac087c2",
  1461 => x"ce059a72",
  1462 => x"c11ec087",
  1463 => x"c049c3dc",
  1464 => x"c487d5f0",
  1465 => x"c087fe86",
  1466 => x"cedcc11e",
  1467 => x"c7f0c049",
  1468 => x"fe1ec087",
  1469 => x"497087e9",
  1470 => x"87fcefc0",
  1471 => x"f887dcc3",
  1472 => x"534f268e",
  1473 => x"61662044",
  1474 => x"64656c69",
  1475 => x"6f42002e",
  1476 => x"6e69746f",
  1477 => x"2e2e2e67",
  1478 => x"e7c01e00",
  1479 => x"f3c087e7",
  1480 => x"87f687cc",
  1481 => x"c21e4f26",
  1482 => x"c048cce8",
  1483 => x"c8e8c278",
  1484 => x"fd78c048",
  1485 => x"87e187fd",
  1486 => x"4f2648c0",
  1487 => x"78452080",
  1488 => x"80007469",
  1489 => x"63614220",
  1490 => x"10df006b",
  1491 => x"2a210000",
  1492 => x"00000000",
  1493 => x"0010df00",
  1494 => x"002a3f00",
  1495 => x"00000000",
  1496 => x"000010df",
  1497 => x"00002a5d",
  1498 => x"df000000",
  1499 => x"7b000010",
  1500 => x"0000002a",
  1501 => x"10df0000",
  1502 => x"2a990000",
  1503 => x"00000000",
  1504 => x"0010df00",
  1505 => x"002ab700",
  1506 => x"00000000",
  1507 => x"000010df",
  1508 => x"00002ad5",
  1509 => x"df000000",
  1510 => x"00000010",
  1511 => x"00000000",
  1512 => x"11740000",
  1513 => x"00000000",
  1514 => x"00000000",
  1515 => x"0017b100",
  1516 => x"4f4f4200",
  1517 => x"20202054",
  1518 => x"4d4f5220",
  1519 => x"616f4c00",
  1520 => x"2e2a2064",
  1521 => x"f0fe1e00",
  1522 => x"cd78c048",
  1523 => x"26097909",
  1524 => x"fe1e1e4f",
  1525 => x"487ebff0",
  1526 => x"1e4f2626",
  1527 => x"c148f0fe",
  1528 => x"1e4f2678",
  1529 => x"c048f0fe",
  1530 => x"1e4f2678",
  1531 => x"52c04a71",
  1532 => x"0e4f2652",
  1533 => x"5d5c5b5e",
  1534 => x"7186f40e",
  1535 => x"7e6d974d",
  1536 => x"974ca5c1",
  1537 => x"a6c8486c",
  1538 => x"c4486e58",
  1539 => x"c505a866",
  1540 => x"c048ff87",
  1541 => x"caff87e6",
  1542 => x"49a5c287",
  1543 => x"714b6c97",
  1544 => x"6b974ba3",
  1545 => x"7e6c974b",
  1546 => x"80c1486e",
  1547 => x"c758a6c8",
  1548 => x"58a6cc98",
  1549 => x"fe7c9770",
  1550 => x"487387e1",
  1551 => x"4d268ef4",
  1552 => x"4b264c26",
  1553 => x"5e0e4f26",
  1554 => x"f40e5c5b",
  1555 => x"d84c7186",
  1556 => x"ffc34a66",
  1557 => x"4ba4c29a",
  1558 => x"73496c97",
  1559 => x"517249a1",
  1560 => x"6e7e6c97",
  1561 => x"c880c148",
  1562 => x"98c758a6",
  1563 => x"7058a6cc",
  1564 => x"ff8ef454",
  1565 => x"1e1e87ca",
  1566 => x"e087e8fd",
  1567 => x"c0494abf",
  1568 => x"0299c0e0",
  1569 => x"1e7287cb",
  1570 => x"49f3ebc2",
  1571 => x"c487f7fe",
  1572 => x"87fdfc86",
  1573 => x"c2fd7e70",
  1574 => x"4f262687",
  1575 => x"f3ebc21e",
  1576 => x"87c7fd49",
  1577 => x"49f6e1c1",
  1578 => x"c487dafc",
  1579 => x"4f2687ff",
  1580 => x"5c5b5e0e",
  1581 => x"ecc20e5d",
  1582 => x"c14abfd2",
  1583 => x"49bfc4e4",
  1584 => x"71bc724c",
  1585 => x"87dbfc4d",
  1586 => x"49744bc0",
  1587 => x"d50299d0",
  1588 => x"d0497587",
  1589 => x"c01e7199",
  1590 => x"fce9c11e",
  1591 => x"1282734a",
  1592 => x"87e4c049",
  1593 => x"2cc186c8",
  1594 => x"abc8832d",
  1595 => x"87daff04",
  1596 => x"c187e8fb",
  1597 => x"c248c4e4",
  1598 => x"78bfd2ec",
  1599 => x"4c264d26",
  1600 => x"4f264b26",
  1601 => x"00000000",
  1602 => x"48d0ff1e",
  1603 => x"ff78e1c8",
  1604 => x"78c548d4",
  1605 => x"c30266c4",
  1606 => x"78e0c387",
  1607 => x"c60266c8",
  1608 => x"48d4ff87",
  1609 => x"ff78f0c3",
  1610 => x"787148d4",
  1611 => x"c848d0ff",
  1612 => x"e0c078e1",
  1613 => x"1e4f2678",
  1614 => x"ebc21e73",
  1615 => x"f2fa49f3",
  1616 => x"c04a7087",
  1617 => x"c204aab7",
  1618 => x"e0c387cd",
  1619 => x"87c905aa",
  1620 => x"48e0e7c1",
  1621 => x"fec178c1",
  1622 => x"aaf0c387",
  1623 => x"c187c905",
  1624 => x"c148dce7",
  1625 => x"87dfc178",
  1626 => x"bfe0e7c1",
  1627 => x"7287c702",
  1628 => x"b3c0c24b",
  1629 => x"4b7287c2",
  1630 => x"bfdce7c1",
  1631 => x"87e0c002",
  1632 => x"b7c44973",
  1633 => x"e8c19129",
  1634 => x"4a7381fc",
  1635 => x"92c29acf",
  1636 => x"307248c1",
  1637 => x"baff4a70",
  1638 => x"98694872",
  1639 => x"87db7970",
  1640 => x"b7c44973",
  1641 => x"e8c19129",
  1642 => x"4a7381fc",
  1643 => x"92c29acf",
  1644 => x"307248c3",
  1645 => x"69484a70",
  1646 => x"c17970b0",
  1647 => x"c048e0e7",
  1648 => x"dce7c178",
  1649 => x"c278c048",
  1650 => x"f849f3eb",
  1651 => x"4a7087e5",
  1652 => x"03aab7c0",
  1653 => x"c087f3fd",
  1654 => x"87e4fc48",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"494a711e",
  1658 => x"2687ccfd",
  1659 => x"4ac01e4f",
  1660 => x"91c44972",
  1661 => x"81fce8c1",
  1662 => x"82c179c0",
  1663 => x"04aab7d0",
  1664 => x"4f2687ee",
  1665 => x"5c5b5e0e",
  1666 => x"4d710e5d",
  1667 => x"7587d4f7",
  1668 => x"2ab7c44a",
  1669 => x"fce8c192",
  1670 => x"cf4c7582",
  1671 => x"6a94c29c",
  1672 => x"2b744b49",
  1673 => x"48c29bc3",
  1674 => x"4c703074",
  1675 => x"4874bcff",
  1676 => x"7a709871",
  1677 => x"7387e4f6",
  1678 => x"87c0fb48",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"25261e16",
  1696 => x"3e3d362e",
  1697 => x"48d0ff1e",
  1698 => x"7178e1c8",
  1699 => x"08d4ff48",
  1700 => x"1e4f2678",
  1701 => x"c848d0ff",
  1702 => x"487178e1",
  1703 => x"7808d4ff",
  1704 => x"ff4866c4",
  1705 => x"267808d4",
  1706 => x"4a711e4f",
  1707 => x"1e4966c4",
  1708 => x"deff4972",
  1709 => x"48d0ff87",
  1710 => x"2678e0c0",
  1711 => x"711e4f26",
  1712 => x"aab7c24a",
  1713 => x"8287c303",
  1714 => x"82ce87c2",
  1715 => x"721e66c4",
  1716 => x"87d5ff49",
  1717 => x"1e4f2626",
  1718 => x"c34ad4ff",
  1719 => x"d0ff7aff",
  1720 => x"78e1c848",
  1721 => x"ebc27ade",
  1722 => x"497abffd",
  1723 => x"7028c848",
  1724 => x"d048717a",
  1725 => x"717a7028",
  1726 => x"7028d848",
  1727 => x"48d0ff7a",
  1728 => x"2678e0c0",
  1729 => x"5b5e0e4f",
  1730 => x"710e5d5c",
  1731 => x"fdebc24c",
  1732 => x"744b4dbf",
  1733 => x"9b66d02b",
  1734 => x"66d483c1",
  1735 => x"87c204ab",
  1736 => x"4a744bc0",
  1737 => x"724966d0",
  1738 => x"75b9ff31",
  1739 => x"72487399",
  1740 => x"484a7030",
  1741 => x"ecc2b071",
  1742 => x"dafe58c1",
  1743 => x"264d2687",
  1744 => x"264b264c",
  1745 => x"d0ff1e4f",
  1746 => x"78c9c848",
  1747 => x"d4ff4871",
  1748 => x"4f267808",
  1749 => x"494a711e",
  1750 => x"d0ff87eb",
  1751 => x"2678c848",
  1752 => x"1e731e4f",
  1753 => x"ecc24b71",
  1754 => x"c302bfcd",
  1755 => x"87ebc287",
  1756 => x"c848d0ff",
  1757 => x"497378c9",
  1758 => x"ffb1e0c0",
  1759 => x"787148d4",
  1760 => x"48c1ecc2",
  1761 => x"66c878c0",
  1762 => x"c387c502",
  1763 => x"87c249ff",
  1764 => x"ecc249c0",
  1765 => x"66cc59c9",
  1766 => x"c587c602",
  1767 => x"c44ad5d5",
  1768 => x"ffffcf87",
  1769 => x"cdecc24a",
  1770 => x"cdecc25a",
  1771 => x"c478c148",
  1772 => x"264d2687",
  1773 => x"264b264c",
  1774 => x"5b5e0e4f",
  1775 => x"710e5d5c",
  1776 => x"c9ecc24a",
  1777 => x"9a724cbf",
  1778 => x"4987cb02",
  1779 => x"edc191c8",
  1780 => x"83714bd7",
  1781 => x"f1c187c4",
  1782 => x"4dc04bd7",
  1783 => x"99744913",
  1784 => x"bfc5ecc2",
  1785 => x"48d4ffb9",
  1786 => x"b7c17871",
  1787 => x"b7c8852c",
  1788 => x"87e804ad",
  1789 => x"bfc1ecc2",
  1790 => x"c280c848",
  1791 => x"fe58c5ec",
  1792 => x"731e87ef",
  1793 => x"134b711e",
  1794 => x"cb029a4a",
  1795 => x"fe497287",
  1796 => x"4a1387e7",
  1797 => x"87f5059a",
  1798 => x"1e87dafe",
  1799 => x"bfc1ecc2",
  1800 => x"c1ecc249",
  1801 => x"78a1c148",
  1802 => x"a9b7c0c4",
  1803 => x"ff87db03",
  1804 => x"ecc248d4",
  1805 => x"c278bfc5",
  1806 => x"49bfc1ec",
  1807 => x"48c1ecc2",
  1808 => x"c478a1c1",
  1809 => x"04a9b7c0",
  1810 => x"d0ff87e5",
  1811 => x"c278c848",
  1812 => x"c048cdec",
  1813 => x"004f2678",
  1814 => x"00000000",
  1815 => x"00000000",
  1816 => x"5f5f0000",
  1817 => x"00000000",
  1818 => x"03000303",
  1819 => x"14000003",
  1820 => x"7f147f7f",
  1821 => x"0000147f",
  1822 => x"6b6b2e24",
  1823 => x"4c00123a",
  1824 => x"6c18366a",
  1825 => x"30003256",
  1826 => x"77594f7e",
  1827 => x"0040683a",
  1828 => x"03070400",
  1829 => x"00000000",
  1830 => x"633e1c00",
  1831 => x"00000041",
  1832 => x"3e634100",
  1833 => x"0800001c",
  1834 => x"1c1c3e2a",
  1835 => x"00082a3e",
  1836 => x"3e3e0808",
  1837 => x"00000808",
  1838 => x"60e08000",
  1839 => x"00000000",
  1840 => x"08080808",
  1841 => x"00000808",
  1842 => x"60600000",
  1843 => x"40000000",
  1844 => x"0c183060",
  1845 => x"00010306",
  1846 => x"4d597f3e",
  1847 => x"00003e7f",
  1848 => x"7f7f0604",
  1849 => x"00000000",
  1850 => x"59716342",
  1851 => x"0000464f",
  1852 => x"49496322",
  1853 => x"1800367f",
  1854 => x"7f13161c",
  1855 => x"0000107f",
  1856 => x"45456727",
  1857 => x"0000397d",
  1858 => x"494b7e3c",
  1859 => x"00003079",
  1860 => x"79710101",
  1861 => x"0000070f",
  1862 => x"49497f36",
  1863 => x"0000367f",
  1864 => x"69494f06",
  1865 => x"00001e3f",
  1866 => x"66660000",
  1867 => x"00000000",
  1868 => x"66e68000",
  1869 => x"00000000",
  1870 => x"14140808",
  1871 => x"00002222",
  1872 => x"14141414",
  1873 => x"00001414",
  1874 => x"14142222",
  1875 => x"00000808",
  1876 => x"59510302",
  1877 => x"3e00060f",
  1878 => x"555d417f",
  1879 => x"00001e1f",
  1880 => x"09097f7e",
  1881 => x"00007e7f",
  1882 => x"49497f7f",
  1883 => x"0000367f",
  1884 => x"41633e1c",
  1885 => x"00004141",
  1886 => x"63417f7f",
  1887 => x"00001c3e",
  1888 => x"49497f7f",
  1889 => x"00004141",
  1890 => x"09097f7f",
  1891 => x"00000101",
  1892 => x"49417f3e",
  1893 => x"00007a7b",
  1894 => x"08087f7f",
  1895 => x"00007f7f",
  1896 => x"7f7f4100",
  1897 => x"00000041",
  1898 => x"40406020",
  1899 => x"7f003f7f",
  1900 => x"361c087f",
  1901 => x"00004163",
  1902 => x"40407f7f",
  1903 => x"7f004040",
  1904 => x"060c067f",
  1905 => x"7f007f7f",
  1906 => x"180c067f",
  1907 => x"00007f7f",
  1908 => x"41417f3e",
  1909 => x"00003e7f",
  1910 => x"09097f7f",
  1911 => x"3e00060f",
  1912 => x"7f61417f",
  1913 => x"0000407e",
  1914 => x"19097f7f",
  1915 => x"0000667f",
  1916 => x"594d6f26",
  1917 => x"0000327b",
  1918 => x"7f7f0101",
  1919 => x"00000101",
  1920 => x"40407f3f",
  1921 => x"00003f7f",
  1922 => x"70703f0f",
  1923 => x"7f000f3f",
  1924 => x"3018307f",
  1925 => x"41007f7f",
  1926 => x"1c1c3663",
  1927 => x"01416336",
  1928 => x"7c7c0603",
  1929 => x"61010306",
  1930 => x"474d5971",
  1931 => x"00004143",
  1932 => x"417f7f00",
  1933 => x"01000041",
  1934 => x"180c0603",
  1935 => x"00406030",
  1936 => x"7f414100",
  1937 => x"0800007f",
  1938 => x"0603060c",
  1939 => x"8000080c",
  1940 => x"80808080",
  1941 => x"00008080",
  1942 => x"07030000",
  1943 => x"00000004",
  1944 => x"54547420",
  1945 => x"0000787c",
  1946 => x"44447f7f",
  1947 => x"0000387c",
  1948 => x"44447c38",
  1949 => x"00000044",
  1950 => x"44447c38",
  1951 => x"00007f7f",
  1952 => x"54547c38",
  1953 => x"0000185c",
  1954 => x"057f7e04",
  1955 => x"00000005",
  1956 => x"a4a4bc18",
  1957 => x"00007cfc",
  1958 => x"04047f7f",
  1959 => x"0000787c",
  1960 => x"7d3d0000",
  1961 => x"00000040",
  1962 => x"fd808080",
  1963 => x"0000007d",
  1964 => x"38107f7f",
  1965 => x"0000446c",
  1966 => x"7f3f0000",
  1967 => x"7c000040",
  1968 => x"0c180c7c",
  1969 => x"0000787c",
  1970 => x"04047c7c",
  1971 => x"0000787c",
  1972 => x"44447c38",
  1973 => x"0000387c",
  1974 => x"2424fcfc",
  1975 => x"0000183c",
  1976 => x"24243c18",
  1977 => x"0000fcfc",
  1978 => x"04047c7c",
  1979 => x"0000080c",
  1980 => x"54545c48",
  1981 => x"00002074",
  1982 => x"447f3f04",
  1983 => x"00000044",
  1984 => x"40407c3c",
  1985 => x"00007c7c",
  1986 => x"60603c1c",
  1987 => x"3c001c3c",
  1988 => x"6030607c",
  1989 => x"44003c7c",
  1990 => x"3810386c",
  1991 => x"0000446c",
  1992 => x"60e0bc1c",
  1993 => x"00001c3c",
  1994 => x"5c746444",
  1995 => x"0000444c",
  1996 => x"773e0808",
  1997 => x"00004141",
  1998 => x"7f7f0000",
  1999 => x"00000000",
  2000 => x"3e774141",
  2001 => x"02000808",
  2002 => x"02030101",
  2003 => x"7f000102",
  2004 => x"7f7f7f7f",
  2005 => x"08007f7f",
  2006 => x"3e1c1c08",
  2007 => x"7f7f7f3e",
  2008 => x"1c3e3e7f",
  2009 => x"0008081c",
  2010 => x"7c7c1810",
  2011 => x"00001018",
  2012 => x"7c7c3010",
  2013 => x"10001030",
  2014 => x"78606030",
  2015 => x"4200061e",
  2016 => x"3c183c66",
  2017 => x"78004266",
  2018 => x"c6c26a38",
  2019 => x"6000386c",
  2020 => x"00600000",
  2021 => x"0e006000",
  2022 => x"5d5c5b5e",
  2023 => x"4c711e0e",
  2024 => x"bfdeecc2",
  2025 => x"c04bc04d",
  2026 => x"02ab741e",
  2027 => x"a6c487c7",
  2028 => x"c578c048",
  2029 => x"48a6c487",
  2030 => x"66c478c1",
  2031 => x"ee49731e",
  2032 => x"86c887df",
  2033 => x"ef49e0c0",
  2034 => x"a5c487ef",
  2035 => x"f0496a4a",
  2036 => x"c6f187f0",
  2037 => x"c185cb87",
  2038 => x"abb7c883",
  2039 => x"87c7ff04",
  2040 => x"264d2626",
  2041 => x"264b264c",
  2042 => x"4a711e4f",
  2043 => x"5ae2ecc2",
  2044 => x"48e2ecc2",
  2045 => x"fe4978c7",
  2046 => x"4f2687dd",
  2047 => x"711e731e",
  2048 => x"aab7c04a",
  2049 => x"c287d303",
  2050 => x"05bfcdcd",
  2051 => x"4bc187c4",
  2052 => x"4bc087c2",
  2053 => x"5bd1cdc2",
  2054 => x"cdc287c4",
  2055 => x"cdc25ad1",
  2056 => x"c14abfcd",
  2057 => x"a2c0c19a",
  2058 => x"87e8ec49",
  2059 => x"cdc248fc",
  2060 => x"fe78bfcd",
  2061 => x"711e87ef",
  2062 => x"1e66c44a",
  2063 => x"fde94972",
  2064 => x"4f262687",
  2065 => x"cdcdc21e",
  2066 => x"d7e649bf",
  2067 => x"d6ecc287",
  2068 => x"78bfe848",
  2069 => x"48d2ecc2",
  2070 => x"c278bfec",
  2071 => x"4abfd6ec",
  2072 => x"99ffc349",
  2073 => x"722ab7c8",
  2074 => x"c2b07148",
  2075 => x"2658deec",
  2076 => x"5b5e0e4f",
  2077 => x"710e5d5c",
  2078 => x"87c8ff4b",
  2079 => x"48d1ecc2",
  2080 => x"497350c0",
  2081 => x"7087fde5",
  2082 => x"9cc24c49",
  2083 => x"cb49eecb",
  2084 => x"497087c3",
  2085 => x"d1ecc24d",
  2086 => x"c105bf97",
  2087 => x"66d087e2",
  2088 => x"daecc249",
  2089 => x"d60599bf",
  2090 => x"4966d487",
  2091 => x"bfd2ecc2",
  2092 => x"87cb0599",
  2093 => x"cbe54973",
  2094 => x"02987087",
  2095 => x"c187c1c1",
  2096 => x"87c0fe4c",
  2097 => x"d8ca4975",
  2098 => x"02987087",
  2099 => x"ecc287c6",
  2100 => x"50c148d1",
  2101 => x"97d1ecc2",
  2102 => x"e3c005bf",
  2103 => x"daecc287",
  2104 => x"66d049bf",
  2105 => x"d6ff0599",
  2106 => x"d2ecc287",
  2107 => x"66d449bf",
  2108 => x"caff0599",
  2109 => x"e4497387",
  2110 => x"987087ca",
  2111 => x"87fffe05",
  2112 => x"dcfb4874",
  2113 => x"5b5e0e87",
  2114 => x"f40e5d5c",
  2115 => x"4c4dc086",
  2116 => x"c47ebfec",
  2117 => x"ecc248a6",
  2118 => x"c178bfde",
  2119 => x"c71ec01e",
  2120 => x"87cdfd49",
  2121 => x"987086c8",
  2122 => x"ff87cd02",
  2123 => x"87ccfb49",
  2124 => x"e349dac1",
  2125 => x"4dc187ce",
  2126 => x"97d1ecc2",
  2127 => x"87c302bf",
  2128 => x"c287fed4",
  2129 => x"4bbfd6ec",
  2130 => x"bfcdcdc2",
  2131 => x"87e9c005",
  2132 => x"e249fdc3",
  2133 => x"fac387ee",
  2134 => x"87e8e249",
  2135 => x"ffc34973",
  2136 => x"c01e7199",
  2137 => x"87cefb49",
  2138 => x"b7c84973",
  2139 => x"c11e7129",
  2140 => x"87c2fb49",
  2141 => x"fac586c8",
  2142 => x"daecc287",
  2143 => x"029b4bbf",
  2144 => x"cdc287dd",
  2145 => x"c749bfc9",
  2146 => x"987087d7",
  2147 => x"c087c405",
  2148 => x"c287d24b",
  2149 => x"fcc649e0",
  2150 => x"cdcdc287",
  2151 => x"c287c658",
  2152 => x"c048c9cd",
  2153 => x"c2497378",
  2154 => x"87cd0599",
  2155 => x"e149ebc3",
  2156 => x"497087d2",
  2157 => x"c20299c2",
  2158 => x"734cfb87",
  2159 => x"0599c149",
  2160 => x"f4c387cd",
  2161 => x"87fce049",
  2162 => x"99c24970",
  2163 => x"fa87c202",
  2164 => x"c849734c",
  2165 => x"87cd0599",
  2166 => x"e049f5c3",
  2167 => x"497087e6",
  2168 => x"d40299c2",
  2169 => x"e2ecc287",
  2170 => x"87c902bf",
  2171 => x"c288c148",
  2172 => x"c258e6ec",
  2173 => x"c14cff87",
  2174 => x"c449734d",
  2175 => x"87ce0599",
  2176 => x"ff49f2c3",
  2177 => x"7087fddf",
  2178 => x"0299c249",
  2179 => x"ecc287db",
  2180 => x"487ebfe2",
  2181 => x"03a8b7c7",
  2182 => x"486e87cb",
  2183 => x"ecc280c1",
  2184 => x"c2c058e6",
  2185 => x"c14cfe87",
  2186 => x"49fdc34d",
  2187 => x"87d4dfff",
  2188 => x"99c24970",
  2189 => x"c287d502",
  2190 => x"02bfe2ec",
  2191 => x"c287c9c0",
  2192 => x"c048e2ec",
  2193 => x"87c2c078",
  2194 => x"4dc14cfd",
  2195 => x"ff49fac3",
  2196 => x"7087f1de",
  2197 => x"0299c249",
  2198 => x"ecc287d9",
  2199 => x"c748bfe2",
  2200 => x"c003a8b7",
  2201 => x"ecc287c9",
  2202 => x"78c748e2",
  2203 => x"fc87c2c0",
  2204 => x"c04dc14c",
  2205 => x"c003acb7",
  2206 => x"66c487d1",
  2207 => x"82d8c14a",
  2208 => x"c6c0026a",
  2209 => x"744b6a87",
  2210 => x"c00f7349",
  2211 => x"1ef0c31e",
  2212 => x"f749dac1",
  2213 => x"86c887db",
  2214 => x"c0029870",
  2215 => x"a6c887e2",
  2216 => x"e2ecc248",
  2217 => x"66c878bf",
  2218 => x"c491cb49",
  2219 => x"80714866",
  2220 => x"bf6e7e70",
  2221 => x"87c8c002",
  2222 => x"c84bbf6e",
  2223 => x"0f734966",
  2224 => x"c0029d75",
  2225 => x"ecc287c8",
  2226 => x"f349bfe2",
  2227 => x"cdc287c9",
  2228 => x"c002bfd1",
  2229 => x"c24987dd",
  2230 => x"987087c7",
  2231 => x"87d3c002",
  2232 => x"bfe2ecc2",
  2233 => x"87eff249",
  2234 => x"cff449c0",
  2235 => x"d1cdc287",
  2236 => x"f478c048",
  2237 => x"87e9f38e",
  2238 => x"5c5b5e0e",
  2239 => x"711e0e5d",
  2240 => x"deecc24c",
  2241 => x"cdc149bf",
  2242 => x"d1c14da1",
  2243 => x"747e6981",
  2244 => x"87cf029c",
  2245 => x"744ba5c4",
  2246 => x"deecc27b",
  2247 => x"c8f349bf",
  2248 => x"747b6e87",
  2249 => x"87c4059c",
  2250 => x"87c24bc0",
  2251 => x"49734bc1",
  2252 => x"d487c9f3",
  2253 => x"87c70266",
  2254 => x"7087da49",
  2255 => x"c087c24a",
  2256 => x"d5cdc24a",
  2257 => x"d8f2265a",
  2258 => x"00000087",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"4a711e00",
  2262 => x"49bfc8ff",
  2263 => x"2648a172",
  2264 => x"c8ff1e4f",
  2265 => x"c0fe89bf",
  2266 => x"c0c0c0c0",
  2267 => x"87c401a9",
  2268 => x"87c24ac0",
  2269 => x"48724ac1",
  2270 => x"5e0e4f26",
  2271 => x"0e5d5c5b",
  2272 => x"d4ff4b71",
  2273 => x"4866d04c",
  2274 => x"49d678c0",
  2275 => x"87f4dbff",
  2276 => x"6c7cffc3",
  2277 => x"99ffc349",
  2278 => x"c3494d71",
  2279 => x"e0c199f0",
  2280 => x"87cb05a9",
  2281 => x"6c7cffc3",
  2282 => x"d098c348",
  2283 => x"c3780866",
  2284 => x"4a6c7cff",
  2285 => x"c331c849",
  2286 => x"4a6c7cff",
  2287 => x"4972b271",
  2288 => x"ffc331c8",
  2289 => x"714a6c7c",
  2290 => x"c84972b2",
  2291 => x"7cffc331",
  2292 => x"b2714a6c",
  2293 => x"c048d0ff",
  2294 => x"9b7378e0",
  2295 => x"7287c202",
  2296 => x"2648757b",
  2297 => x"264c264d",
  2298 => x"1e4f264b",
  2299 => x"5e0e4f26",
  2300 => x"f80e5c5b",
  2301 => x"c81e7686",
  2302 => x"fdfd49a6",
  2303 => x"7086c487",
  2304 => x"c0486e4b",
  2305 => x"c6c301a8",
  2306 => x"c34a7387",
  2307 => x"d0c19af0",
  2308 => x"87c702aa",
  2309 => x"05aae0c1",
  2310 => x"7387f4c2",
  2311 => x"0299c849",
  2312 => x"c6ff87c3",
  2313 => x"c34c7387",
  2314 => x"05acc29c",
  2315 => x"c487cdc1",
  2316 => x"31c94966",
  2317 => x"66c41e71",
  2318 => x"c292d44a",
  2319 => x"7249e6ec",
  2320 => x"e0d5fe81",
  2321 => x"4966c487",
  2322 => x"49e3c01e",
  2323 => x"87d9d9ff",
  2324 => x"d8ff49d8",
  2325 => x"c0c887ee",
  2326 => x"d6dbc21e",
  2327 => x"f5f1fd49",
  2328 => x"48d0ff87",
  2329 => x"c278e0c0",
  2330 => x"d01ed6db",
  2331 => x"92d44a66",
  2332 => x"49e6ecc2",
  2333 => x"d3fe8172",
  2334 => x"86d087e8",
  2335 => x"c105acc1",
  2336 => x"66c487cd",
  2337 => x"7131c949",
  2338 => x"4a66c41e",
  2339 => x"ecc292d4",
  2340 => x"817249e6",
  2341 => x"87cdd4fe",
  2342 => x"1ed6dbc2",
  2343 => x"d44a66c8",
  2344 => x"e6ecc292",
  2345 => x"fe817249",
  2346 => x"c887f4d1",
  2347 => x"c01e4966",
  2348 => x"d7ff49e3",
  2349 => x"49d787f3",
  2350 => x"87c8d7ff",
  2351 => x"c21ec0c8",
  2352 => x"fd49d6db",
  2353 => x"d087feef",
  2354 => x"48d0ff86",
  2355 => x"f878e0c0",
  2356 => x"87d1fc8e",
  2357 => x"5c5b5e0e",
  2358 => x"711e0e5d",
  2359 => x"4cd4ff4d",
  2360 => x"487e66d4",
  2361 => x"06a8b7c3",
  2362 => x"48c087c5",
  2363 => x"7587e2c1",
  2364 => x"c1e2fe49",
  2365 => x"c41e7587",
  2366 => x"93d44b66",
  2367 => x"83e6ecc2",
  2368 => x"ccfe4973",
  2369 => x"83c887fd",
  2370 => x"d0ff4b6b",
  2371 => x"78e1c848",
  2372 => x"49737cdd",
  2373 => x"7199ffc3",
  2374 => x"c849737c",
  2375 => x"ffc329b7",
  2376 => x"737c7199",
  2377 => x"29b7d049",
  2378 => x"7199ffc3",
  2379 => x"d849737c",
  2380 => x"7c7129b7",
  2381 => x"7c7c7cc0",
  2382 => x"7c7c7c7c",
  2383 => x"7c7c7c7c",
  2384 => x"78e0c07c",
  2385 => x"dc1e66c4",
  2386 => x"dcd5ff49",
  2387 => x"7386c887",
  2388 => x"cefa2648",
  2389 => x"5b5e0e87",
  2390 => x"1e0e5d5c",
  2391 => x"d4ff7e71",
  2392 => x"c21e6e4b",
  2393 => x"fe49faec",
  2394 => x"c487d8cb",
  2395 => x"9d4d7086",
  2396 => x"87c3c302",
  2397 => x"bfc2edc2",
  2398 => x"fe496e4c",
  2399 => x"ff87f7df",
  2400 => x"c5c848d0",
  2401 => x"7bd6c178",
  2402 => x"7b154ac0",
  2403 => x"e0c082c1",
  2404 => x"f504aab7",
  2405 => x"48d0ff87",
  2406 => x"c5c878c4",
  2407 => x"7bd3c178",
  2408 => x"78c47bc1",
  2409 => x"c1029c74",
  2410 => x"dbc287fc",
  2411 => x"c0c87ed6",
  2412 => x"b7c08c4d",
  2413 => x"87c603ac",
  2414 => x"4da4c0c8",
  2415 => x"e8c24cc0",
  2416 => x"49bf97c7",
  2417 => x"d20299d0",
  2418 => x"c21ec087",
  2419 => x"fe49faec",
  2420 => x"c487cccd",
  2421 => x"4a497086",
  2422 => x"c287efc0",
  2423 => x"c21ed6db",
  2424 => x"fe49faec",
  2425 => x"c487f8cc",
  2426 => x"4a497086",
  2427 => x"c848d0ff",
  2428 => x"d4c178c5",
  2429 => x"bf976e7b",
  2430 => x"c1486e7b",
  2431 => x"c17e7080",
  2432 => x"f0ff058d",
  2433 => x"48d0ff87",
  2434 => x"9a7278c4",
  2435 => x"c087c505",
  2436 => x"87e5c048",
  2437 => x"ecc21ec1",
  2438 => x"cafe49fa",
  2439 => x"86c487e0",
  2440 => x"fe059c74",
  2441 => x"d0ff87c4",
  2442 => x"78c5c848",
  2443 => x"c07bd3c1",
  2444 => x"c178c47b",
  2445 => x"c087c248",
  2446 => x"4d262648",
  2447 => x"4b264c26",
  2448 => x"5e0e4f26",
  2449 => x"710e5c5b",
  2450 => x"0266cc4b",
  2451 => x"c04c87d8",
  2452 => x"d8028cf0",
  2453 => x"c14a7487",
  2454 => x"87d1028a",
  2455 => x"87cd028a",
  2456 => x"87c9028a",
  2457 => x"497387d7",
  2458 => x"d087eafb",
  2459 => x"c01e7487",
  2460 => x"87e0f949",
  2461 => x"49731e74",
  2462 => x"c887d9f9",
  2463 => x"87fcfe86",
  2464 => x"dac21e00",
  2465 => x"c149bfea",
  2466 => x"eedac2b9",
  2467 => x"48d4ff59",
  2468 => x"ff78ffc3",
  2469 => x"e1c848d0",
  2470 => x"48d4ff78",
  2471 => x"31c478c1",
  2472 => x"d0ff7871",
  2473 => x"78e0c048",
  2474 => x"00004f26",
  2475 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
